XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I�@W�(�n�r�1�&br�
F.~�`\�u>���NՏ��>&�3Q�q�1@R���u����q>�o�������q���2�&�%�q��v���*R���*��7*
�7�L����������{ �9�rlؑ�4���PI�3�50xaQ�lp��E�ɬYn�K#?�yhK&+2a�Q�
��o�a:+x��R
l�)Y�}ג��������t}i� 
1$�6�g��$��N�	M��u�Y�w�[��H���a���c����Y�_G���<��	�nJx��{���2��2�e$�1ƭ�@�\Luf�A2^M�il���cC۪�L�u�B��oq����^���+��=�4�l����z�r�{�7��a�3���������~�(#�*���c���
D>�S
/�����Qn�*ǖ��B76pÏ��+�.�;?a[_g�O�4D8��ݼ���U�l�Nb�EM}Z�s+b$̼\�b���68��CS��("�©���-�&�q'��H}D������k@�VBʜ�����M6�v�<���s�k��J���&���74�B�\����@?v�����7�,��
���I3M�Ic(�G2�F���?$��X*��͜һx^5��nT���,��;Oa'��T����x���$�u�N�pl��K��m"�1)Cc<r��^K6]�?!�����*�wG�7�,w�U�f��90���;$��b����_�`�x���V"b^�r�Y�N�d�BYכ�XlxVHYEB    1602     7a0�%�\pg����z��JA)KiB��f_��ˎD�pyg(�n庳t1F��͢1��FZCIH(���>��X'��͸���	��!�:Q066�@��x �����&�֯A{��U�N7�����-:�[�[	���{���g���'�3v]]�5�o�����"�U��o6aT �_�}��q7?�3��x
|3��'����[>�c/����}\Cm:����HN�OE��Hb�Q��\|PH�z���a�����
�G�}�t����IVD��	�N�{�N!1�T�IP��}�|	�[����/W��tf<c�v��K����8w9�ga��iY�J���,��[����*Ř��������i�"`C��&Y0y�q�k�.π1ة|9t[yK._� ʐ��C��é�ڈ����U�[�C�}/g�����#�o���<�i���;�.�(���FuO��Vt��c�
�e���I۶�E�Z�d�𷴍F���5����ib�d�j�T	"�<������0"����!��6��Aw�[bl�R=>��?�5�L�M�ӷD^��Y�%:$(�گo16�M�c��d�gCOҡpa����pO^�wYes�����s�f�Ƨ�p������X��J]�㩝l�Y�"]�Fc����`P�j��\��5�_E�Md��8�of\H^�E�����F�c^��z_�V�D����u�g�p���?w��ѯ�F�Y#����Q�!j�,����Nu���t���%&�	;t����^�_k��ƛ]7 ����0*<+��>`��$����Q���5X��y���:	{w��$I.F��� �I��7Ke��[�njũ=�)��p��"�f�O�`]�4zaYm'�I���t��}yg#aݵ�F8D͟�/d1�9��Cл]��$#*޿~?�ѥꁮ��Y^n�k5��i�6�����^Q@�/,��R��.��WCe�3���q�x��j�DGC��H���^�ʩn*�d2�p>����x�6(�D	�9��$.� 5���6��u��c�b*3�i�=��~�H�U�!��ŪS���A'*�BuN���ol��u���N����BP�;�[�8���+Έ���I�.���b7.	jYb�J��C����LƑ������[�	�M�щ��`�o�h��Gt&<KT�����h*	�7�]�(�/J
hs0�4���J�f+����e��C�QA�E�����ŗ��Ӧ;X�J�3K$q�����b��ʊZ�q�i��$�d%��`�}J�J�xv��;��L[n�+��˴�����v�Ğwr���*��w^y����H�|���5�uŠ�
n��u˖��&���%Q.��wky��u��V,z�#+,�(ޡ���Lc��Y�@�Z>�ԫ���pK!� .I��ޙ��[�jA@���~HD�(sm����E�e��s�:�y��)��~l�����!�c�i5�����0�g��`L��]�A�ѷ¾d����ޖCGN�$�ۃJaSz�-e|�-���Ď���G�T����]j� �������\l��r�6r�'(����$FȜ%�kp�֜�bJ�����Q�O|�0�%l1Zå�3�C7��r�텫k�Fi�:K�.�(=Cqr4��66�b䟻��XMeT�c�(n�k?����>X��!��li�v ��c�rc ]�rQ+H��{���T4s�ζ;����[�>n054�@.P��"�Z⎦1��4�ǗE�!�,��c#�� �y��{�.q��{g����� #���j�������x���+�� �)���I���E߱����Ҋ�B%x9_�(�<����sK����Ծn�������L8�8F��������?��ej7���Ձ�`Q�ז���ƈ�&