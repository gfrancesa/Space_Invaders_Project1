XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���G�($5�
%�mņ��@c�r��[j���=���O�a���7�V�;���:�Q4�'_�n�~���|�,�MǸ^O3���d�S��?Y�Ԥ7/���s����F�yg����:ý�J5�C�Z�Np:�9zPpQ��i5�ƿyv&���xt|��|4�ʻ8q+��L�{�h�`�Y�H��P`����~� �P�Ў�r����*����A��q��5���Y�����y�`&[ 7?E�y씱\V"�'t7��}��ɏ"�v�{��W@(���.+;�7 �Yc4�{���o����k�e#�n�7$�����a�#�[�4e$R�{�(^2$vm��f��ձ���~q@:ü�Z����7Hj6����@.�*R%[��Ԭ;�)�k���(I�2������R�"++�{
z:�\�_��B�� ��u�����:jZ�@ĵr�!u�Y�S�69�.����Fo�o��T�ώr���i��X%��g�ln-�<(�"�v z�J�r�hT�����e��8y�D7V�Y��ac��Z�3kvpMݯwm��3r�b"���̞�I����=�Cs�𛣙�db1eE%�sX��8��Y���녻[D��+��K�|���kϨ)_s� �|�V�t-x��@��CO�d[A����1�7��b'�`9���+�ˎ�*֭�(+�6]=��hp2���A�-z�ʋ�b2(��?j|�K7���#���z7�/G���ӭH�7��,���È�f�nV��ph���XlxVHYEB    3189     890��������ŧ�Y���u�g�ˌs��05�V[�\��+O ��"צ�V�Tk������e������:[޼ۂ4�?�����wL�ӁT_o욶F���Dq�������k�B�-`*��\�sN�Wp2���q�Ze��C�.mOL3�Еe0kKM�u����"ҳiV${	j�;��Lc@U����D��.|�Ww��F��^�m�>g	��v�FX� l�7�!�r�յ��Y�2�Y׫7�S�w��FTd/��,�8=�0&�k73Y����;�_ͥ#':.A�maM%�(�q+���߆W�'�\�M��_�=���՘9WB�W6���u���Q�(C�~�67a~Y��1�P@`���#�J������r�9�tL\V|%��q��KZ'l��㧤�Ս.��:��N�����dPb:�Ε������C�����-0F�oi1�Ѯ��.����o���𘺚	!���G�<�N�.��Bt�L�85(m!�+愚X��*�hCe�LG���9����R͂�u�b�#O�B�Y����)��= �	Hn���9��.]ف��n�����\�W��ID�^&�a�J:���/���>O�G�ܓ�p�a����+�q?��t�D���j�n˙Qޜ�߄��Щ/�3C��U�u
��&v�Q�E&S�`���a��D��1��|�����+�t>��,���m-	x��sbo9 ���9T�k����R��v�y�
{�<�s�T�ߍXn̕qs�������0�����/�c`ezC%ۮ<��}�@��b��̮��SlHaƀ�#E
9��'� �����&��n��j������m���^��Nѧ~ ��&I	B9��r�s���Q���@Nkz��}�(I��6ersLU�K��(�b?��4�cٍ,Ir-fԹ���&����'�("��x�1���ǖ���E�Θ�#f(bu�x}$�a��2Է ��U����+��Gu���B��LT��)��E~����nA�[e�P,� _�eD>��@����D?bvy���@H�T`��ݚ���� ͔Q:$6z0
��E��ħ��٩�%�>u��--��ö����_�̔[^�U�|�����^a:8-���,$՞�GG6�?�n�E�{�!�e˗s.X��Z��jg�[�ϚWkeg�n� ��)��(4���>)�ؼ=ׅ��M�6k���:ߝ���訄Ȅ�ݤ�7�|������:���z�����V�C�$�_	�e�D��S��1���""��V��fM�}M*�Y�D���{%[������"�CEp�#��{�8�I�dj!i����^��4�4;G��)�鎁�>�jS��Q�2�e��E�Wz��3~!�>�%������Vj�G�1�d�8�8������vN�l�*��&{��S��5�|!~� ,�`����`�¶+�PV�tI�P��<l�б����<�Z����4��Fi��(q�ڷ����~�O�"o|E�C���eT�_�r�db0�)�ۀi�_�eEC�ݗhSJ�r��G���p�۷͙fM	V�c9p�!�m@-a��]D�zr�S�;�7�o�Nh�.?��Z���W���Z�{qi#G��`W9U.o�>����[�U!$z=�)K^�c�{�.�#��wp7st�6���H��.�<!�wD����sG֥$�n�t�+��p����=�賦�s��F`>L�^��`g8R8��q��>_�	V��֙�N�F�;=d�|w斢Ү��2����������t��j�4�(�&��z�3#�=�Im�����Ģ�jEw3t���c2|P+���ܱ[k��۠AM;�λ����_���N�+T3W8��~9��*�Y����ރo3�������*f�_�P�١Y��T<���"�2���*	�j�����݄/C�`i�Yϋh@{��c��+����a�x� ����J�jTfH�8{�\4���4M���zkx��t&��ICd2����R����Jbݐ^
Bޚ Ӝ�H�(k'JdduK	4?2]�i�ү��S.���Ѻ^ƅ�0L�fu2�(U��i-���e�.��	�e�7At��VķU5/��"Z�\���5?����iq���m� ���o5��	9D]@�.3r