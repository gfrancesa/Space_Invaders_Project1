`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:56:26 10/26/2014 
// Design Name: 
// Module Name:    Figures_ROM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Figures_ROM(
			input wire clk,
			input wire [10:0] addr,
			output reg [31:0] data
    );
   
   // signal declaration
   reg [10:0] addr_reg; 

   // body
   always @(posedge clk) 
      addr_reg <= addr;
      
   always @*
      case (addr_reg)
         //code x00
			
			11'h000: data = 32'b00000000000000000000000000000000; // 
         11'h001: data = 32'b00000000000000000000000000000000; // 
         11'h002: data = 32'b00000000000000000000000000000000; //   ****
         11'h003: data = 32'b00000000000000000000000000000000; //  **  **
         11'h004: data = 32'b00000000000000000000000000000000; //  **  **
         11'h005: data = 32'b00000000000000000000000000000000; //  **  **
         11'h006: data = 32'b00000000000000000000000000000000; //  **  **
         11'h007: data = 32'b00000000000000111100000000000000; //   ****
         11'h008: data = 32'b00000000000000111100000000000000; //    **
         11'h009: data = 32'b00000000000011111111000000000000; //  ******
         11'h00a: data = 32'b00000000000011111111000000000000; //    **
         11'h00b: data = 32'b00000000001111111111110000000000; //    **
         11'h00c: data = 32'b00000000001111111111110000000000; // 
         11'h00d: data = 32'b00000000111100111100111100000000; // 
         11'h00e: data = 32'b00000000111100111100111100000000; // 
         11'h00f: data = 32'b00000000111111111111111100000000; // 
         11'h010: data = 32'b00000000111111111111111100000000; // 
         11'h011: data = 32'b00000000000011000011000000000000; // 
         11'h012: data = 32'b00000000000011000011000000000000; //   ******
         11'h013: data = 32'b00000000001100111100110000000000; //   **  **
         11'h014: data = 32'b00000000001100111100110000000000; //   ******
         11'h015: data = 32'b00000000110011000011001100000000; //   **
         11'h016: data = 32'b00000000110011000011001100000000; //   **
         11'h017: data = 32'b00000000000000000000000000000000; //   **
         11'h018: data = 32'b00000000000000000000000000000000; //   **
         11'h019: data = 32'b00000000000000000000000000000000; //  ***
         11'h01a: data = 32'b00000000000000000000000000000000; // ****
         11'h01b: data = 32'b00000000000000000000000000000000; // ***
         11'h01c: data = 32'b00000000000000000000000000000000; // 
         11'h01d: data = 32'b00000000000000000000000000000000; // 
         11'h01e: data = 32'b00000000000000000000000000000000; // 
         11'h01f: data = 32'b00000000000000000000000000000000; //
			// ------------------------------------------------------------------------------

         //code x07
         11'h020: data = 32'b00000000000000000000000000000000; // 
         11'h021: data = 32'b00000000000000000000000000000000; // 
         11'h022: data = 32'b00000000000000000000000000000000; //  *******
         11'h023: data = 32'b00000000000000000000000000000000; //  **   **
         11'h024: data = 32'b00000000000000000000000000000000; //  *******
         11'h025: data = 32'b00000000000000000000000000000000; //  **   **
         11'h026: data = 32'b00000000000000000000000000000000; //  **   **
         11'h027: data = 32'b00000000011000000000011000000000; //  **   **////
         11'h028: data = 32'b00000000011000000000011000000000; //  **   **
         11'h029: data = 32'b00000110000110000001100001100000; //  **  ***
         11'h02a: data = 32'b00000110000110000001100001100000; // ***  ***
         11'h02b: data = 32'b00000110011111111111111001100000; // ***  **
         11'h02c: data = 32'b00000110011111111111111001100000; // **
         11'h02d: data = 32'b00000111111001111110011111100000; // 
         11'h02e: data = 32'b00000111111001111110011111100000; // 
         11'h02f: data = 32'b00000111111111111111111111100000; // 
         11'h030: data = 32'b00000111111111111111111111100000; // 
         11'h031: data = 32'b00000001111111111111111110000000; // 
         11'h032: data = 32'b00000001111111111111111110000000; // 
         11'h033: data = 32'b00000000011000000000011000000000; //    **
         11'h034: data = 32'b00000000011000000000011000000000; //    **
         11'h035: data = 32'b00000001100000000000000110000000; // ** ** **
         11'h036: data = 32'b00000001100000000000000110000000; //   ****
         11'h037: data = 32'b00000000000000000000000000000000; // ***  ***
         11'h038: data = 32'b00000000000000000000000000000000; //   ****
         11'h039: data = 32'b00000000000000000000000000000000; // ** ** **
         11'h03a: data = 32'b00000000000000000000000000000000; //    **
         11'h03b: data = 32'b00000000000000000000000000000000; //    **
         11'h03c: data = 32'b00000000000000000000000000000000; // 
         11'h03d: data = 32'b00000000000000000000000000000000; // 
         11'h03e: data = 32'b00000000000000000000000000000000; // 
         11'h03f: data = 32'b00000000000000000000000000000000; // 
         //code x08
         11'h040: data = 32'b00000000000000000000000000000000; // 
         11'h041: data = 32'b00000000000000000000000000000000; // *
         11'h042: data = 32'b00000000000000000000000000000000; // **
         11'h043: data = 32'b00000000000000000000000000000000; // ***
         11'h044: data = 32'b00000000000000000000000000000000; // ****
         11'h045: data = 32'b00000000000000000000000000000000; // *****
         11'h046: data = 32'b00000000000000000000000000000000; // *******
         11'h047: data = 32'b00000000000000000000000000000000; // ***** 
         11'h048: data = 32'b00000000000011111111000000000000; // **** //
         11'h049: data = 32'b00000000000011111111000000000000; // ***
         11'h04a: data = 32'b00000011111111111111111111000000; // **
         11'h04b: data = 32'b00000011111111111111111111000000; // *
         11'h04c: data = 32'b00001111111111111111111111110000; // 
         11'h04d: data = 32'b00001111111111111111111111110000; // 
         11'h04e: data = 32'b00001111110000111100001111110000; // 
         11'h04f: data = 32'b00001111110000111100001111110000; // 
         11'h050: data = 32'b00001111111111111111111111110000; // 
         11'h051: data = 32'b00001111111111111111111111110000; //       *
         11'h052: data = 32'b00000000001111000011110000000000; //      **
         11'h053: data = 32'b00000000001111000011110000000000; //     ***
         11'h054: data = 32'b00000000111100111100111100000000; //    ****
         11'h055: data = 32'b00000000111100111100111100000000; //   *****
         11'h056: data = 32'b00001111000000000000000011110000; // *******
         11'h057: data = 32'b00001111000000000000000011110000; //   *****
         11'h058: data = 32'b00000000000000000000000000000000; //    ****
         11'h059: data = 32'b00000000000000000000000000000000; //     ***
         11'h05a: data = 32'b00000000000000000000000000000000; //      **
         11'h05b: data = 32'b00000000000000000000000000000000; //       *
         11'h05c: data = 32'b00000000000000000000000000000000; // 
         11'h05d: data = 32'b00000000000000000000000000000000; // 
         11'h05e: data = 32'b00000000000000000000000000000000; // 
         11'h05f: data = 32'b00000000000000000000000000000000; // 





			// -------------------------------------------------------------------------------
			 
			 
			 
			 
			 
			 
			 
			 
			 
			 
			11'h060: data = 32'b00000000000000000000000000000000; // 
         11'h061: data = 32'b00000000000000000000000000000000; // 
         11'h062: data = 32'b00000000000000000000000000000000; //    **
         11'h063: data = 32'b00000000000000000000000000000000; //   ****
         11'h064: data = 32'b00000000000000000000000000000000; //  ******
         11'h065: data = 32'b00000000000000000000000000000000; //    **
         11'h066: data = 32'b00000000000000000000000000000000; //    **
         11'h067: data = 32'b00000000000000000000000000000000; //    **
         11'h068: data = 32'b00000000000000000000000000000000; //    **
         11'h069: data = 32'b00000000000000000000000000000000; //    **
         11'h06a: data = 32'b00000000000000110000000000000000; //    **
         11'h06b: data = 32'b00000000000000110000000000000000; //    **
         11'h06c: data = 32'b00000000000011111100000000000000; // 
         11'h06d: data = 32'b00000000000011111100000000000000; // 
         11'h06e: data = 32'b00001111111111111111111111110000; // 
         11'h06f: data = 32'b00001111111111111111111111110000; // 
         11'h070: data = 32'b00111111111111111111111111111100; // 
         11'h071: data = 32'b00111111111111111111111111111100; // 
         11'h072: data = 32'b00111111111111111111111111111100; //    **
         11'h073: data = 32'b00111111111111111111111111111100; //    **
         11'h074: data = 32'b00111111111111111111111111111100; //    **
         11'h075: data = 32'b00111111111111111111111111111100; //    **
         11'h076: data = 32'b00111111111111111111111111111100; //    **
         11'h077: data = 32'b00111111111111111111111111111100; //    **
         11'h078: data = 32'b00000000000000000000000000000000; //    **
         11'h079: data = 32'b00000000000000000000000000000000; //  ******
         11'h07a: data = 32'b00000000000000000000000000000000; //   ****
         11'h07b: data = 32'b00000000000000000000000000000000; //    **
         11'h07c: data = 32'b00000000000000000000000000000000; // 
         11'h07d: data = 32'b00000000000000000000000000000000; // 
         11'h07e: data = 32'b00000000000000000000000000000000; // 
         11'h07f: data = 32'b00000000000000000000000000000000; // 
 
         //code x04
         11'h080: data = 32'b00000000000000000000000000000000; // ********
         11'h081: data = 32'b00000000000000000000000000000000; // ********
         11'h082: data = 32'b00000000000000000000000000000000; // ********
         11'h083: data = 32'b00000000000000000000000000000000; // ********
         11'h084: data = 32'b00000000000000000000000000000000; // ********
         11'h085: data = 32'b00000000000000000000000000000000; // ********
         11'h086: data = 32'b00000000000000000000000000000000; // ***  ***
         11'h087: data = 32'b00000000000000000000000000000000; // **    **
         11'h088: data = 32'b00000000000000000000000000000000; // **    **
         11'h089: data = 32'b00000000000000000000000000000000; // ***  ***
         11'h08a: data = 32'b00000000000000000000000000000000; // ********
         11'h08b: data = 32'b00000000000000000000000000000000; // ********
         11'h08c: data = 32'b00000000000000000000000000000000; // ********
         11'h08d: data = 32'b00000000000000000000000000000000; // ********
         11'h08e: data = 32'b00000000000000000000000000000000; // ********
         11'h08f: data = 32'b00000000000000000000000000000000; // ********
         11'h090: data = 32'b00000000000000000000000000000000; // 
         11'h091: data = 32'b00000000000000000000000000000000; // 
         11'h092: data = 32'b00000000000000000000000000000000; // 
         11'h093: data = 32'b00000000000000000000000000000000; // 
         11'h094: data = 32'b00000000000000000000000000000000; // 
         11'h095: data = 32'b00000000000000000000000000000000; //   ****
         11'h096: data = 32'b00000000000000000000000000000000; //  **  **
         11'h097: data = 32'b00000000000000000000000000000000; //  *    *
         11'h098: data = 32'b00000000000000000000000000000000; //  *    *
         11'h099: data = 32'b00000000000000000000000000000000; //  **  **
         11'h09a: data = 32'b00000000000000000000000000000000; //   ****
         11'h09b: data = 32'b00000000000000000000000000000000; // 
         11'h09c: data = 32'b00000000000000000000000000000000; // 
         11'h09d: data = 32'b00000000000000000000000000000000; // 
         11'h09e: data = 32'b00000000000000000000000000000000; // 
         11'h09f: data = 32'b00000000000000000000000000000000; // 
         //code x05
         11'h0a0: data = 32'b00000000000000000000000000001111; // ********
         11'h0a1: data = 32'b00000000000000000000000000001111; // ********
         11'h0a2: data = 32'b00000000000000000000000000001111; // ********
         11'h0a3: data = 32'b00000000000000000000000000001111; // ********
         11'h0a4: data = 32'b00000000000000000000000000001111; // ********
         11'h0a5: data = 32'b00000000000000000000000000001111; // **    **
         11'h0a6: data = 32'b00000000000000000000000000001111; // *  **  *
         11'h0a7: data = 32'b00000000000000000000000000001111; // * **** *
         11'h0a8: data = 32'b00000000000000000000000000001111; // * **** *
         11'h0a9: data = 32'b00000000000000000000000000001111; // *  **  *
         11'h0aa: data = 32'b00000000000000000000000000001111; // **    **
         11'h0ab: data = 32'b00000000000000000000000000001111; // ********
         11'h0ac: data = 32'b00000000000000000000000000001111; // ********
         11'h0ad: data = 32'b00000000000000000000000000001111; // ********
         11'h0ae: data = 32'b00000000000000000000000000001111; // ********
         11'h0af: data = 32'b00000000000000000000000000001111; // ********
         11'h0b0: data = 32'b00000000000000000000000000001111; // 
         11'h0b1: data = 32'b00000000000000000000000000001111; // 
         11'h0b2: data = 32'b00000000000000000000000000001111; //    ****
         11'h0b3: data = 32'b00000000000000000000000000001111; //     ***
         11'h0b4: data = 32'b00000000000000000000000000001111; //    ** *
         11'h0b5: data = 32'b00000000000000000000000000001111; //   **  *
         11'h0b6: data = 32'b00000000000000000000000000001111; //  ****
         11'h0b7: data = 32'b00000000000000000000000000001111; // **  **
         11'h0b8: data = 32'b00000000000000000000000000001111; // **  **
         11'h0b9: data = 32'b00000000000000000000000000001111; // **  **
         11'h0ba: data = 32'b00000000000000000000000000001111; // **  **
         11'h0bb: data = 32'b00000000000000000000000000001111; //  ****
         11'h0bc: data = 32'b00000000000000000000000000001111; // 
         11'h0bd: data = 32'b00000000000000000000000000001111; // 
         11'h0be: data = 32'b00000000000000000000000000001111; // 
         11'h0bf: data = 32'b00000000000000000000000000001111; // 
         //code x06
         11'h0c0: data = 32'b00000000000011111111000000000000; // 
         11'h0c1: data = 32'b00000000000011111111000000000000; // 
         11'h0c2: data = 32'b00000000000011111111000000000000; //   ****
         11'h0c3: data = 32'b00000000000011111111000000000000; //  **  **
         11'h0c4: data = 32'b00000000111111111111111100000000; //  **  **
         11'h0c5: data = 32'b00000000111111111111111100000000; //  **  **
         11'h0c6: data = 32'b00000000111111111111111100000000; //  **  **
         11'h0c7: data = 32'b00000000111111111111111100000000; //   ****
         11'h0c8: data = 32'b00001111111111111111111111110000; //    **
         11'h0c9: data = 32'b00001111111111111111111111110000; //  ******
         11'h0ca: data = 32'b00001111111111111111111111110000; //    **
         11'h0cb: data = 32'b00001111111111111111111111110000; //    **
         11'h0cc: data = 32'b11111111000011111111000011111111; // 
         11'h0cd: data = 32'b11111111000011111111000011111111; // 
         11'h0ce: data = 32'b11111111000011111111000011111111; // 
         11'h0cf: data = 32'b11111111000011111111000011111111; // 
         11'h0d0: data = 32'b11111111111111111111111111111111; // 
         11'h0d1: data = 32'b11111111111111111111111111111111; // 
         11'h0d2: data = 32'b11111111111111111111111111111111; //   ******
         11'h0d3: data = 32'b11111111111111111111111111111111; //   **  **
         11'h0d4: data = 32'b00000000111100000000111100000000; //   ******
         11'h0d5: data = 32'b00000000111100000000111100000000; //   **
         11'h0d6: data = 32'b00000000111100000000111100000000; //   **
         11'h0d7: data = 32'b00000000111100000000111100000000; //   **
         11'h0d8: data = 32'b00001111000011111111000011110000; //   **
         11'h0d9: data = 32'b00001111000011111111000011110000; //  ***
         11'h0da: data = 32'b00001111000011111111000011110000; // ****
         11'h0db: data = 32'b00001111000011111111000011110000; // ***
         11'h0dc: data = 32'b11110000111100000000111100001111; // 
         11'h0dd: data = 32'b11110000111100000000111100001111; // 
         11'h0de: data = 32'b11110000111100000000111100001111; // 
         11'h0df: data = 32'b11110000111100000000111100001111; // 
         //code x07
         11'h0e0: data = 32'b00000000000000000000000000000000; // 
         11'h0e1: data = 32'b00000000000000000000000000000000; // 
         11'h0e2: data = 32'b00000000000000000000000000000000; //  *******
         11'h0e3: data = 32'b00000000000000000000000000000000; //  **   **
         11'h0e4: data = 32'b00000000000000000000000000000000; //  *******
         11'h0e5: data = 32'b00000000000000000000000000000000; //  **   **
         11'h0e6: data = 32'b00000000000000000000000000000000; //  **   **
         11'h0e7: data = 32'b00000000011000000000011000000000; //  **   **////
         11'h0e8: data = 32'b00000000011000000000011000000000; //  **   **
         11'h0e9: data = 32'b00000110000110000001100001100000; //  **  ***
         11'h0ea: data = 32'b00000110000110000001100001100000; // ***  ***
         11'h0eb: data = 32'b00000110011111111111111001100000; // ***  **
         11'h0ec: data = 32'b00000110011111111111111001100000; // **
         11'h0ed: data = 32'b00000111111001111110011111100000; // 
         11'h0ee: data = 32'b00000111111001111110011111100000; // 
         11'h0ef: data = 32'b00000111111111111111111111100000; // 
         11'h0f0: data = 32'b00000111111111111111111111100000; // 
         11'h0f1: data = 32'b00000001111111111111111110000000; // 
         11'h0f2: data = 32'b00000001111111111111111110000000; // 
         11'h0f3: data = 32'b00000000011000000000011000000000; //    **
         11'h0f4: data = 32'b00000000011000000000011000000000; //    **
         11'h0f5: data = 32'b00000001100000000000000110000000; // ** ** **
         11'h0f6: data = 32'b00000001100000000000000110000000; //   ****
         11'h0f7: data = 32'b00000000000000000000000000000000; // ***  ***
         11'h0f8: data = 32'b00000000000000000000000000000000; //   ****
         11'h0f9: data = 32'b00000000000000000000000000000000; // ** ** **
         11'h0fa: data = 32'b00000000000000000000000000000000; //    **
         11'h0fb: data = 32'b00000000000000000000000000000000; //    **
         11'h0fc: data = 32'b00000000000000000000000000000000; // 
         11'h0fd: data = 32'b00000000000000000000000000000000; // 
         11'h0fe: data = 32'b00000000000000000000000000000000; // 
         11'h0ff: data = 32'b00000000000000000000000000000000; // 
         //code x08
         11'h100: data = 32'b00000000000000000000000000000000; // 
         11'h101: data = 32'b00000000000000000000000000000000; // *
         11'h102: data = 32'b00000000000000000000000000000000; // **
         11'h103: data = 32'b00000000000000000000000000000000; // ***
         11'h104: data = 32'b00000000000000000000000000000000; // ****
         11'h105: data = 32'b00000000000000000000000000000000; // *****
         11'h106: data = 32'b00000000000000000000000000000000; // *******
         11'h107: data = 32'b00000000000000000000000000000000; // ***** 
         11'h108: data = 32'b00000000000011111111000000000000; // **** //
         11'h109: data = 32'b00000000000011111111000000000000; // ***
         11'h10a: data = 32'b00000011111111111111111111000000; // **
         11'h10b: data = 32'b00000011111111111111111111000000; // *
         11'h10c: data = 32'b00001111111111111111111111110000; // 
         11'h10d: data = 32'b00001111111111111111111111110000; // 
         11'h10e: data = 32'b00001111110000111100001111110000; // 
         11'h10f: data = 32'b00001111110000111100001111110000; // 
         11'h110: data = 32'b00001111111111111111111111110000; // 
         11'h111: data = 32'b00001111111111111111111111110000; //       *
         11'h112: data = 32'b00000000001111000011110000000000; //      **
         11'h113: data = 32'b00000000001111000011110000000000; //     ***
         11'h114: data = 32'b00000000111100111100111100000000; //    ****
         11'h115: data = 32'b00000000111100111100111100000000; //   *****
         11'h116: data = 32'b00001111000000000000000011110000; // *******
         11'h117: data = 32'b00001111000000000000000011110000; //   *****
         11'h118: data = 32'b00000000000000000000000000000000; //    ****
         11'h119: data = 32'b00000000000000000000000000000000; //     ***
         11'h11a: data = 32'b00000000000000000000000000000000; //      **
         11'h11b: data = 32'b00000000000000000000000000000000; //       *
         11'h11c: data = 32'b00000000000000000000000000000000; // 
         11'h11d: data = 32'b00000000000000000000000000000000; // 
         11'h11e: data = 32'b00000000000000000000000000000000; // 
         11'h11f: data = 32'b00000000000000000000000000000000; // 
         //code x09
         11'h120: data = 32'b00000000000011111111000000000000; // 
         11'h121: data = 32'b00000000000011111111000000000000; // 
         11'h122: data = 32'b00000000000011111111000000000000; //    **
         11'h123: data = 32'b00000000000011111111000000000000; //   ****
         11'h124: data = 32'b00000000111111111111111100000000; //  ******
         11'h125: data = 32'b00000000111111111111111100000000; //    **
         11'h126: data = 32'b00000000111111111111111100000000; //    **
         11'h127: data = 32'b00000000111111111111111100000000; //    **
         11'h128: data = 32'b00001111111111111111111111110000; //  ******
         11'h129: data = 32'b00001111111111111111111111110000; //   ****
         11'h12a: data = 32'b00001111111111111111111111110000; //    **
         11'h12b: data = 32'b00001111111111111111111111110000; // 
         11'h12c: data = 32'b11111111000011111111000011111111; // 
         11'h12d: data = 32'b11111111000011111111000011111111; // 
         11'h12e: data = 32'b11111111000011111111000011111111; // 
         11'h12f: data = 32'b11111111000011111111000011111111; // 
         11'h130: data = 32'b11111111111111111111111111111111; // 
         11'h131: data = 32'b11111111111111111111111111111111; // 
         11'h132: data = 32'b11111111111111111111111111111111; //  **  **
         11'h133: data = 32'b11111111111111111111111111111111; //  **  **
         11'h134: data = 32'b00001111000011111111000011110000; //  **  **
         11'h135: data = 32'b00001111000011111111000011110000; //  **  **
         11'h136: data = 32'b00001111000011111111000011110000; //  **  **
         11'h137: data = 32'b00001111000011111111000011110000; //  **  **
         11'h138: data = 32'b11110000000000000000000000001111; //  **  **
         11'h139: data = 32'b11110000000000000000000000001111; // 
         11'h13a: data = 32'b11110000000000000000000000001111; //  **  **
         11'h13b: data = 32'b11110000000000000000000000001111; //  **  **
         11'h13c: data = 32'b00001111000000000000000011110000; // 
         11'h13d: data = 32'b00001111000000000000000011110000; // 
         11'h13e: data = 32'b00001111000000000000000011110000; // 
         11'h13f: data = 32'b00001111000000000000000011110000; // 
         //code x10
         11'h140: data = 32'b00000000000000000000000000000000; // 
         11'h141: data = 32'b00000000000000000000000000000000; // 
         11'h142: data = 32'b00000000000000000000000000000000; //  *******
         11'h143: data = 32'b00000000000000000000000000000000; // ** ** **
         11'h144: data = 32'b00000000000000000000000000000000; // ** ** **
         11'h145: data = 32'b00000000000000000000000000000000; // ** ** **
         11'h146: data = 32'b00000000000000000000000000000000; //  **** **
         11'h147: data = 32'b00000000000000000000000000000000; //    ** **
         11'h148: data = 32'b00000000011000000000011000000000; //    ** **
         11'h149: data = 32'b00000000011000000000011000000000; //    ** **
         11'h14a: data = 32'b00000000000110000001100000000000; //    ** **
         11'h14b: data = 32'b00000000000110000001100000000000; //    ** **
         11'h14c: data = 32'b00000000011111111111111000000000; // 
         11'h14d: data = 32'b00000000011111111111111000000000; // 
         11'h14e: data = 32'b00000001111001111110011110000000; // 
         11'h14f: data = 32'b00000001111001111110011110000000; // 
         11'h150: data = 32'b00000111111111111111111111100000; // 
         11'h151: data = 32'b00000111111111111111111111100000; //  *****
         11'h152: data = 32'b00000110011111111111111001100000; // **   **
         11'h153: data = 32'b00000110011111111111111001100000; //  **
         11'h154: data = 32'b00000110011000000000001101100000; //   ***
         11'h155: data = 32'b00000110011000000000001101100000; //  ** **
         11'h156: data = 32'b00000000000111100011110000000000; // **   **
         11'h157: data = 32'b00000000000111100011110000000000; // **   **
         11'h158: data = 32'b00000000000000000000000000000000; //  ** **
         11'h159: data = 32'b00000000000000000000000000000000; //   ***
         11'h15a: data = 32'b00000000000000000000000000000000; //     **
         11'h15b: data = 32'b00000000000000000000000000000000; // **   **
         11'h15c: data = 32'b00000000000000000000000000000000; //  *****
         11'h15d: data = 32'b00000000000000000000000000000000; // 
         11'h15e: data = 32'b00000000000000000000000000000000; // 
         11'h15f: data = 32'b00000000000000000000000000000000; // 
         //code x11
         11'h160: data = 32'b00000000000000000000000000000000; // 
         11'h161: data = 32'b00000000000000000000000000000000; // 
         11'h162: data = 32'b00000000000000000000000000000000; // 
         11'h163: data = 32'b00000000000000000000000000000000; // 
         11'h164: data = 32'b00000000000000000000000000000000; // 
         11'h165: data = 32'b00000000000000000000000000000000; // 
         11'h166: data = 32'b00000000000000000000000000000000; // 
         11'h167: data = 32'b00000000000000000000000000000000; // 
         11'h168: data = 32'b00000000000011111111000000000000; // *******
         11'h169: data = 32'b00000000000011111111000000000000; // *******
         11'h16a: data = 32'b00000011111111111111111111000000; // *******
         11'h16b: data = 32'b00000011111111111111111111000000; // *******
         11'h16c: data = 32'b00001111111111111111111111110000; // 
         11'h16d: data = 32'b00001111111111111111111111110000; // 
         11'h16e: data = 32'b00001111110000111100001111110000; // 
         11'h16f: data = 32'b00001111110000111100001111110000; // 
         11'h170: data = 32'b00001111111111111111111111110000; // 
         11'h171: data = 32'b00001111111111111111111111110000; // 
         11'h172: data = 32'b00000000111111000011111100000000; //    **
         11'h173: data = 32'b00000000111111000011111100000000; //   ****
         11'h174: data = 32'b00000011110000111100001111000000; //  ******
         11'h175: data = 32'b00000011110000111100001111000000; //    **
         11'h176: data = 32'b00000000111100000000111100000000; //    **
         11'h177: data = 32'b00000000111100000000111100000000; //    **
         11'h178: data = 32'b00000000000000000000000000000000; //  ******
         11'h179: data = 32'b00000000000000000000000000000000; //   ****
         11'h17a: data = 32'b00000000000000000000000000000000; //    **
         11'h17b: data = 32'b00000000000000000000000000000000; //  ******
         11'h17c: data = 32'b00000000000000000000000000000000; // 
         11'h17d: data = 32'b00000000000000000000000000000000; // 
         11'h17e: data = 32'b00000000000000000000000000000000; // 
         11'h17f: data = 32'b00000000000000000000000000000000; // 
         //code x12
         11'h180: data = 32'b00000000000000000000000000000000; // 
         11'h181: data = 32'b00000000000000000000000000000000; // 
         11'h182: data = 32'b00000000000000000000000000000000; //    **
         11'h183: data = 32'b00000000000000000000000000000000; //   ****
         11'h184: data = 32'b00000000000000000000000000000000; //  ******
         11'h185: data = 32'b00000000000000000000000000000000; //    **
         11'h186: data = 32'b00000000000000000000000000000000; //    **
         11'h187: data = 32'b00000000000000000000000000000000; //    **
         11'h188: data = 32'b00000000000000000000000000000000; //    **
         11'h189: data = 32'b00000000000000000000000000000000; //    **
         11'h18a: data = 32'b00000000000000110000000000000000; //    **
         11'h18b: data = 32'b00000000000000110000000000000000; //    **
         11'h18c: data = 32'b00000000000011111100000000000000; // 
         11'h18d: data = 32'b00000000000011111100000000000000; // 
         11'h18e: data = 32'b00001111111111111111111111110000; // 
         11'h18f: data = 32'b00001111111111111111111111110000; // 
         11'h190: data = 32'b00111111111111111111111111111100; // 
         11'h191: data = 32'b00111111111111111111111111111100; // 
         11'h192: data = 32'b00111111111111111111111111111100; //    **
         11'h193: data = 32'b00111111111111111111111111111100; //    **
         11'h194: data = 32'b00111111111111111111111111111100; //    **
         11'h195: data = 32'b00111111111111111111111111111100; //    **
         11'h196: data = 32'b00111111111111111111111111111100; //    **
         11'h197: data = 32'b00111111111111111111111111111100; //    **
         11'h198: data = 32'b00000000000000000000000000000000; //    **
         11'h199: data = 32'b00000000000000000000000000000000; //  ******
         11'h19a: data = 32'b00000000000000000000000000000000; //   ****
         11'h19b: data = 32'b00000000000000000000000000000000; //    **
         11'h19c: data = 32'b00000000000000000000000000000000; // 
         11'h19d: data = 32'b00000000000000000000000000000000; // 
         11'h19e: data = 32'b00000000000000000000000000000000; // 
         11'h19f: data = 32'b00000000000000000000000000000000; // 
         //code x13
         11'h1a0: data = 32'b00000000000000000000000000000000; // 
         11'h1a1: data = 32'b00000000000000000000000000000000; // 
         11'h1a2: data = 32'b00000000000000000000000000000000; // 
         11'h1a3: data = 32'b00000000000000000000000000000000; // 
         11'h1a4: data = 32'b00000000000000000000000000000000; // 
         11'h1a5: data = 32'b00000000000000000000000000000000; //    **
         11'h1a6: data = 32'b00000000000000000000000000000000; //     **
         11'h1a7: data = 32'b00000000000000000000000000000000; // *******
         11'h1a8: data = 32'b00000000001111111111110000000000; //     **//
         11'h1a9: data = 32'b00000000001111111111110000000000; //    **
         11'h1aa: data = 32'b00000011111111111111111111000000; // 
         11'h1ab: data = 32'b00000011111111111111111111000000; // 
         11'h1ac: data = 32'b00001111111111111111111111110000; // 
         11'h1ad: data = 32'b00001111111111111111111111110000; // 
         11'h1ae: data = 32'b00111100111100111100111100111100; // 
         11'h1af: data = 32'b00111100111100111100111100111100; // 
         11'h1b0: data = 32'b11111111111111111111111111111111; // 
         11'h1b1: data = 32'b11111111111111111111111111111111; // 
         11'h1b2: data = 32'b00001111110000111100001111110000; // 
         11'h1b3: data = 32'b00001111110000111100001111110000; // 
         11'h1b4: data = 32'b00000011000000000000000011000000; // 
         11'h1b5: data = 32'b00000011000000000000000011000000; //   **
         11'h1b6: data = 32'b00000000000000000000000000000000; //  **
         11'h1b7: data = 32'b00000000000000000000000000000000; // *******
         11'h1b8: data = 32'b00000000000000000000000000000000; //  **
         11'h1b9: data = 32'b00000000000000000000000000000000; //   **
         11'h1ba: data = 32'b00000000000000000000000000000000; // 
         11'h1bb: data = 32'b00000000000000000000000000000000; // 
         11'h1bc: data = 32'b00000000000000000000000000000000; // 
         11'h1bd: data = 32'b00000000000000000000000000000000; // 
         11'h1be: data = 32'b00000000000000000000000000000000; // 
         11'h1bf: data = 32'b00000000000000000000000000000000; // 
         //code x14
         11'h1c0: data = 32'b10000000000000000000000000000000; // 
         11'h1c1: data = 32'b01000000000000000000000000000000; // 
         11'h1c2: data = 32'b00100000000000000000000000000000; // 
         11'h1c3: data = 32'b00010000000000000000000000000000; // 
         11'h1c4: data = 32'b00001000000000000000000000000000; // 
         11'h1c5: data = 32'b00000100000000000000000000000000; // 
         11'h1c6: data = 32'b00000010000000000000000000000000; // **
         11'h1c7: data = 32'b00000001000000000000000000000000; // **
         11'h1c8: data = 32'b00000000100000000000000000000000; // **
         11'h1c9: data = 32'b00000000010000000000000000000000; // *******
         11'h1ca: data = 32'b00000000001000000000000000000000; // 
         11'h1cb: data = 32'b00000000000100000000000000000000; // 
         11'h1cc: data = 32'b00000000000010000000000000000000; // 
         11'h1cd: data = 32'b00000000000001000000000000000000; // 
         11'h1ce: data = 32'b00000000000000100000000000000000; // 
         11'h1cf: data = 32'b00000000000000010000000000000000; // 
         11'h1d0: data = 32'b00000000000000001000000000000000; // 
         11'h1d1: data = 32'b00000000000000000100000000000000; // 
         11'h1d2: data = 32'b00000000000000000010000000000000; // 
         11'h1d3: data = 32'b00000000000000000001000000000000; // 
         11'h1d4: data = 32'b00000000000000000000100000000000; // 
         11'h1d5: data = 32'b00000000000000000000010000000000; //   *  *
         11'h1d6: data = 32'b00000000000000000000001000000000; //  **  **
         11'h1d7: data = 32'b00000000000000000000000100000000; // ********
         11'h1d8: data = 32'b00000000000000000000000010000000; //  **  **
         11'h1d9: data = 32'b00000000000000000000000001000000; //   *  *
         11'h1da: data = 32'b00000000000000000000000000100000; // 
         11'h1db: data = 32'b00000000000000000000000000010000; // 
         11'h1dc: data = 32'b00000000000000000000000000001000; // 
         11'h1dd: data = 32'b00000000000000000000000000000100; // 
         11'h1de: data = 32'b00000000000000000000000000000010; // 
         11'h1df: data = 32'b00000000000000000000000000000001; // 
         //code x15
         11'h1e0: data = 32'b00000000000001000000000000000000; // 
         11'h1e1: data = 32'b00000000000001000000000000000000; // 
         11'h1e2: data = 32'b00000000000001000000000000000000; // 
         11'h1e3: data = 32'b00000000000001000000000000000000; // 
         11'h1e4: data = 32'b00000000000001000000000000000000; //    *
         11'h1e5: data = 32'b00000000000001000000000000000000; //   ***
         11'h1e6: data = 32'b00000000000001000000000000000000; //   ***
         11'h1e7: data = 32'b00000000000001000000000000000000; //  *****
         11'h1e8: data = 32'b00000000000001000000000000000000; //  *****
         11'h1e9: data = 32'b00000000000001000000000000000000; // *******
         11'h1ea: data = 32'b00000000000001000000000000000000; // *******
         11'h1eb: data = 32'b00000000000001000000000000000000; // 
         11'h1ec: data = 32'b00000000000001000000000000000000; // 
         11'h1ed: data = 32'b00000000000001000000000000000000; // 
         11'h1ee: data = 32'b00000000000001000000000000000000; // 
         11'h1ef: data = 32'b00000000000001000000000000000000; // 
         11'h1f0: data = 32'b00000000000001000000000000000000; // 
         11'h1f1: data = 32'b00000000000001000000000000000000; // 
         11'h1f2: data = 32'b00000000000001000000000000000000; // 
         11'h1f3: data = 32'b00000000000001000000000000000000; // 
         11'h1f4: data = 32'b00000000000001000000000000000000; // *******
         11'h1f5: data = 32'b00000000000001000000000000000000; // *******
         11'h1f6: data = 32'b00000000000001000000000000000000; //  *****
         11'h1f7: data = 32'b00000000000001000000000000000000; //  *****
         11'h1f8: data = 32'b00000000000001000000000000000000; //   ***
         11'h1f9: data = 32'b00000000000001000000000000000000; //   ***
         11'h1fa: data = 32'b00000000000001000000000000000000; //    *
         11'h1fb: data = 32'b00000000000001000000000000000000; // 
         11'h1fc: data = 32'b00000000000001000000000000000000; // 
         11'h1fd: data = 32'b00000000000001000000000000000000; // 
         11'h1fe: data = 32'b00000000000001000000000000000000; // 
         11'h1ff: data = 32'b00000000000001000000000000000000; // 
        
        
   	 
   endcase  
   	       
endmodule
