XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����u��qC#�j��j#��ȿ�K!!jS�T,��'�x�bgf��p�N��\���g
�Eȷ�:H�38�2g5m�,�}���od��TO���2k�/���L�ZLq�d3@�u�Q�Ȅ�'������s'A�1��
V,�\D(�q#��.����<�	��2�����)}����m$gv ~�@�ލ��J��n�:�}�sv$���ĩ<��&�80Ы��	HgW��8���w��J����������r-�o^N��{	_�bq$�.4ǹA �8orj������&ת��M7�\0��𵳤_x�SԳy�B��'	�	n>:R���*�����ވ �!-�;��ѐ�܀���o^\T��<�p��E�H��#\�Ԁ
��b���m��2#�a��i�h��u[�G�	��֪E����CDi�y#�A���V�\���<4͙#�{ꬹyF���(Q��4�����NhR�f���rt`�e蚛���F���q~w��I����F� �INי�y�0?�Zz��X�&j����_���y�B\?*�V�����>���n.z:
��G���Ύ�= N�.�|>~0UO�� �Y��"�C`��V����ݥ���6�8�"IJ+�����:Z�@��+�t7�o�Z�q��(g�I���@�xv^�R?׺�1�9������AL�Ac'8!�S���l���7�9QA�]"}W����f���-	Y�NP������YӃ�֋,;�_�|u+FMn rK�XlxVHYEB    3357     c80�cu�Hm=X,�Ux�������'L��;�tH�FU�zS�4��X��ղ���W��єE��MC��&�?�cJ�VJ�k�#h?TF�;��&,(��rf�E��Z���O(�D�L^'@�:k���3g4�f�����B���Է�)���V"�S؎V���aq#��X�];(�
i����i�7kSy���Q̤���K��H§㠲�w�^�o*_��A��8���E�&����<�V"������z y���w|U�g.AGV�[ a�����ǘ�۫mt<V�jχJ_��	��I����[�c\H�@����-#M(���2m.���0�pu/��8s���?E�~K}�W�m7PZ��
9�~�����c�������q��/H�֐! }A�D��#R��%���T�����w��+_4��Qogei_�f��@^�B�U��x���/�Ͳ��~�$.�h2ѠC�@�~wp�X��߉��l\����~[�\�[��}?9��F�	t�����6w�C*	#�ݹO�^�'X�Q`���GL״�Id*@��h����;@F��_�"YPv_ZN����D����&�`��$�q�UY�5�܎����d ���z����6z˟Ȭ�o�:�~�Ӧn�G$p��ΗG�����R���~�l���f�s1l�֡2T�.=�������'�����{͵��=oc����핟1��Ff#ne���%C�a���g9��xߘA����#ҽ,w �/�b�v�F%�$���EP�g ^��~O�R�S�P�}��Q�2a��Z�|�llG�H���F*t��~.v�"��4$���9��Lp�Hf�� �|&�֭*v4P���ި�C��N��Q�V�>�����{��L�=v����u;4���� �~K��#����?���Z��E�F/��yD�� �/�a�*����ۃ+a�gm�1`/���L�c��^߷o�g��@w�'��)��݉�D�B]A��v����7����B�9��`&�}"���9v�b���
�Vҥ��ltpQh���±Q��i�Q���8r�
��n�%���-@���)P����a���q��@�,�T�@�v�,���Jt��g	o�0>�_�C�Zv��2�����
����c!�
�qF��`ryE�k}���*Λ幕�L�����gu�#"Ʌ��1�K�x��w��D����c�!o<�GM V�'�B�������
����nU����|>]-I�>~��"\~v�z��-f����U1�mO5�:ZC>�L�����O�~�>㘯؏Y���u��L3�b��K�E�/����$�2f�w����n��8q�$z{yP���D
;�0�n��*ѝ\��&Md�}kk��f�j�0�#pqԂ{�Y�y�~6�o�<���e*��źLި�SS��m!���}/rV����>Уδ��GN�H�"��������b�Q���͔M��xm��N��;y�s�G7+/�8\�'� �H�Er���f�:�{ ���]p1~p|/HO�E��W��%��H��P)�u(ax)�ḒJ���ʃ��)�d ��Oo��Y(��8~���c�b�΄��^_����g�{3"T�F���Z}�
����*=�B���El5�^�6��.���ʥ2<2�:��%U'Y�+�h+A��0�_{3ޤ?�jF4���~�K�3R`U=����1����3���q�c��>៥��Rd�!T�6�����h�@���J7���އd]�f�0-y�C���iu/�#�ꉀ���_)���^�e���j]ddmB=�Z� 5��4!D�	*s}kׇ�*5Z�!�9��W|1/��P�/�>0��i�"����x�������j�N5"�dj��o�C\S�\�v%�j+-;*M�{�V���Ϧ1, wZ���yi�������m����4���}ӕ�-#��;�_���JS�D���q�Xf�CP���=����9a ��l?Ku��'"'`2z'�� ���X�^��������p�썝�?3;v���T#E$w����d����g���4�|
�=륀��S�V_L�����1]�;g6��j=N5��M��N_gc�|�0ߛk��W��(�F�Ã@3� �<��D��`���k���nș�_��O��)���e��}�N�h�1��J���b�ܽ�u#�V��pz#�9'�*0
�������8 #Zǚ�4N��ԋMc�Fp&�B��t21U����N�襈�sv�f�;R��[�
J4��VY��[�k��Ǥ/�����L:�떝jP�A���&��nA�>H���Lȃ:�g_��7���<]��s�j��Mi�[̩�^��+V
_S���O_%� �}�[�@,!�z?���F�k�*C��3!KCK���n�Mp5�i��Ṍ�$��q~ �ب/J#��G�K%"���F�Y5��:�*�D���	����E�Ɉ�y��N��?֓ۗ��r�$m*�����b�%�^��8OyM=֥΀�;��Z�&�������v��澾��̇(�	��ڨ�o�6'�k���K����%��:]�e��&�7d5Z�M�ꚹ���$e3,��t}v���1���~�EbKo_�'���-jQ���u��D��Q��;�@'��e9YE���D;n��u���[Bu̦�V_����A�T�-��o�H�(���u�b��؁�r!���ַ�=V��8�wOj�͖Xzz��S�%nf�j�mLO�g�a���!����L���i���?[��兓5)�T��u�j4�O'�o]k�IY�`�9�&�-�Ҟġ<�����|�Wřg� |;�;sz�h� uӯW&�g�x�:3��J�c��^la^Ju7�Ix��8u�������%��Ck�v�oH�B����w��� �\����ӏ1�a��7��(��hb&E�_���ȡ��$;Xjf��]�F�z	c�G�A3���/Ķ�������se�(0�`)�d��~�	9:�Trd��	���MjE� �G%+��Z{+Gx��@Tu��d�n��Z�k�gf�&P��?4S&6���܋ą�6�\-Q�C,���{T��eY�튵£T굱��..���>-@3S�'Ҵ���