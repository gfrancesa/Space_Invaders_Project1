XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��wi�G5A;ᴉ9� �1[n��)��k����X�J���3\)|�c@}cÜ�4��\`�m��̖z#�X�b�KFc�ڑ��B��}��yx����2��G.���W<{��1��1�e>��R�e�lB�_�/G3o���*�?�R}s4��ڑa��V6ݒ�-o��@�=�p{P���e�ʏ�i��j]穘c�����?�1�N���]X�C��o��S&>�"!��Xl��8��.�hј��N�5��Z��G)�_�.�̿_��㾰�+Ĝ��}�aħ�	e�˪��f���P����Ll�z�k�I�)h��س���oC�`N��Rz�ڃ5��MK��.x .i~K�	'a�(�b����B�0; (�꽸�Mg��ʀd/�x�
H�=��豷�N0��u��=�!��ޅ����݋�5	3	�+��N�|����J�	�/�I�UwRZH�=cTe8����ڶ۽��$��Q>Ք I��f�b����<��(�l���%�.J��'>�Y�6s�@L��z��<�k�<B��@�Z&��G��t3Vk�H�����0�~PH�xv�"4�=�yQ0-��5�8�R^W��5e�Ӏny��bz�IY��j\�z�3��&���}Q��s��ſ������N�^Èm��gl*mR�]@&`�Gl`J����}aŹb����T���_�0�����)�+��u����Yܥ�u��,w��[%@�^*��fX�/FJw�w�>'�<a:tV=
��׃�6^�XlxVHYEB    5ee8    14d0�ʑ��L&Gyj*˩�G���V��V���s���6��	�����'e24��z(�'�g��X?N�E%_�B�ȭ.�L�ZS�Z�ޱͬRx��c+�-Y)k�	�V~rv�[^���~@(~V�����3 B�mR{\�+�s\�H���l8� =B�{TL�s#
�|E�q�r�[3['?�2�H�=�n6��V%މ��1���M���D9�s�Q�+�g�/R+�cT�sϋ�?�{��+a=��Ew<���L���Ǳ�k���*�������a~�X���1/AR�0R���d�*{���_@%9��P�?��sDL�l�g{�9Rppn0$�`��g�5��"�l
*SK�8p׌}M�t��q3ѡ6	�Cֵ!)�R)� ��I�0�����D+�������A�\��c8e '�� AaFF�(T�\"-<ht매����{	�#)(����u������̓�����K}Y�iX�"7�d��!d��U���1����6�Wb�V���1Sa:<H���%������^��)����nT��uu�eބ�z�OE˻y���h����|f�鼑*�u2�߃�Z�է8&���1�y(̙n�7�������]΂Ҭ�&�e$����������d@0tm@�0�nA��/:x4����R]�v^�K�/�2��F��tj ���.�I�e��'�`�) aov��M��9�#G���*v�/�K�*5F�yg��F�ˆ�e���t�p�/�d	��-�5�ݍZ'�4��4���2bˠ�/n�эȾ������7��N���{%�ߏr_/�@�������k��&V��f?\$[���������
$�·Q�\���(���Ȝ
�j���ŏ���B�Y"P^�KriJ����Q�lkp�p߻����.9��/Mg�fS:��������J ���2�{�g��ߚ����p�]곻��R�R f���	{ݞ�y����o߭����
�v�-Jٸ���7P��}Ao�݅��0G�'F��|J16�{��̽�l�@���� �3����+F�#y�p�5u��*�i��~C�?R�����{6W�����7�L�;KһԺD�G���Vry��d�&���w@�Ww��԰r�����b
b��ٹw`�7�9_=}輦���~�� 8���O�o���[�^SO��(�)e-w���$i�̏���mG��#+�y�I�Hךǀ�׈��˒�8E1�oArls>�����0�l9-|Х�j�{�˸����[s���W����Q�0�4.���d�F�����$��"г �B2����z+�7eBc-��ݺFM�W�#<6��6k�AG|	5�WRw�b�%^	�s)Ϩ���C��].ܱ�3q"[��Ɓ���)FNJ��?�&~4<�D��p-(c�b�k��$M:0 #��m�����o0\�ؗ���b��/�J��N1߉iFV}��[/�f���8�^�����L���2`��٥f"̮r�X�+��łL^����y��,R���Wf.���L���.�y �P���L@�*m��xZ�I�l�ŝ/�������s/|��4F����	g����i�6A3w��d�j�Y���՟kM#��L9�OƸ/����ߚp5�����a]!~�bH��=�{����-ܷ���z���JŇ��Ņ\g� /l��zg@>�Z���1���x<���I3<%LWkq�8�5�g�m="6�?��P�R�igy#B��r?�$�z\�y�t��,?�c�sgk���̕��;^9�=���H:�t�)�.!V��j���I���zD��	}|F8�����V�驅�j�#����A��x�cd�WئV��{�/�%��Q�
����A�E»�H�&A���'"A���\%���s����|���X*3�m�+'�ʮ��GC�7�#_��<�0-g�ђ�y3v�]���F��R�,����?�o,��b^!�O���+pK���;��	/�Bf�en�nr����mR���Z
Z�e���_�[,��{C�Ǐ�z)�]�^q�����(Oh�&q�X�*]�1�7���V>�+�v���ʥNlcB�\�s�-n
s��L��$6�����	a@�@��!Ʊ=N_,{E)_�^q��\a�s|���BK"�� �����j�2p}�)K*�d��>:RQ;�͆���߼\r�)��<�1�Z��	��K\y*�C�അ^�\w�O�v�>��	]gW�M�~�&��@^�zl�~�^D�O�N�Q��]���*>���bo#�O���׍;k�7bʙS�2R�g �&��#�S9g87*N��!<z��LA��#&(�7�AҖ�"즀I)���#
'����ϣ�����YL�����6�JJ�hl|�	^���\��a��o�c}�f���v}|���j/����
�W�V�͓�_5e���2��K y$�Wc�7�H�.�߃�Ƕ�%���jX�3�1�(B��UP�R�U�:�X�SJ�"�ֲjȯ��<��I�W�Y�X�W�
�����@#�O�D��>�%�B8�T)[ZB�g�\�?��Y�{���3��_�
|nY�2�zMܢ�Q��P~���tҴ�	����B@@�%fȅT�+~�JS{n��*z��V+�«*r%�?�]��y�[[�C�����aH��ʶ�N�:߫RMe�vv��Hc,�zΓx�n9Xtp�ڼ����(+E�^��~|��
*�;�x�8a�=����vJ(�E֤ A�b>�k!�_�qf>?�T�T���T��֕-�ns��M�6��]�H]V�\k��c��d��qr�ƒ�6�1���?��;��� e%�^���f����wj">T��S�ZT����/^�ƾ�Tl��QL_gM;A8OG�T/���$�dt��Ν�,�`B�?�;	�P�%�p�I}����m��/��'s�t�aC�?^����M�`\/8%�H9�<�3Y�Uk1u��<��wH�q*Ʃ�.�+�[�Y��n[='xu��Q�o�lp�i9X&��Hp?�6>a��߷�lcO݊Ӵb0���u�A�hE6=�:�q�\ƒ�a�R����{p���J��|���o}��%�ot��_9��\W̪}���ֽd�����0���\�6S!�L�zP�gk7@F8d�t�Ȯ�h��/ō ݩ)K������֌M�.2e��B��*]������d�$��L{�}";��Oz|�b5И_�!W:��o�k����ibǮ6��L.�y&1�g�C��� ~������e�|�ި�~�YCkܑ�V�����-�	x�(q��#���z�$�U��=��M��V�g�]A��tF'��a�������8Y�:�D�QATl�z���s;.26m����Z�芸�v^wZ�nݬ�h��f�U���;�Č^8�����9뢳��K�}N��3�[��PR���t^�����a��r��q;�j��=�ԚUb�N�y���ω9� ^k	�5���l��R@���P�X�?-�#po �<��� ""����ܾ����A��b&Y����#�d��5�OFĢ`��7Ad�����E�Y2������b��
'@T�y�u����p	���)e��{�k���Ї��xѱ�=8��G��w0���pDJR2�zJx���rn�Z��6�
=�J�])s�E�$P����3X�\�1���c͙��L�-��� `�G�x�T�$�un���ƞ7��6�o�jԔ�`wR������8(��ы֪�89o��RȂpS��q�&!%��r�/���;�S�~��E{7�����x#�����.")N�=�0F��çڒ4�8�O0=e�V�iC��9��a�R�(+Q'���T5�>F��Z��P�:�T��#�#�	Z�����&ֆ P�m���B�k��"wޝe���N^s�k3ӫ�@��>� ��(�-���m9,3W�^}K�f���Sa� �続�Er�����K,�x�۔̈�'����E�Ut�k�������N-�°,u=xh�~UEVEF{�,�-9Fc�|�D^�Dr�G�s�3�a��p&^����A�\����p�d-c\���ęa�iqI*p4Uy�^ �ga�h8��zt! ���8��=S���@��_�����2ƺS��k�lt�F�~�6Ҍ��}
�␬_�.T���,��z� ���;i�C��k���@��%���3N�z�-R��uP��=^��8���4�dg�;E��#NT�����O�rO�c뀶>��9K���i�}�[}��؇Xj�W3��p7���(�z�Y.ū�7Zr&B��~j�@��8]��.N���	U<ݪ�(�運Y�_x�(��/u�9+n��'
q�_.�z�9�f��O·<���q�^ߟ����Ds�a�"M�B^���aHʌ��YFi[�$p��N'�����k���E����MC�\o�(H�̿B���� Yʹ��}�Je�ҡ3�k#έ�1��u��4�Ψ_�>�_�ib��4�?D�ɟ����Ή���w�+T��C+0EK�ݹ>���3�愶�#dX�H�x��ZD���� ~�H��`.��]�䗛&pY��Y�BH��l���^V��P����~����A{�l&(��2-ȍh�bj$?qusޔ�f#�D�T�ܗ<NH"��݊]�ET�aQ��o�0�zed���}��v]�oE����$�x�P�n���Y�WCe�n��2��G��hB��4R���W�$�a��wk��܀�^�""��W� ��w)]_�S���� ��F4�+KL� դgoP�u��p҂�"���آr]�A"X���M18V�X���9�7��׀+�+��BvS��)���{X�x
~޷lP��'���uR β�\JV,�nϝD�#Sd���b��~@Y0����2~�2�_IԿ$��O)�.�I���}�F�qU�GH~gV���(�A��¾��9�b.�d���P��6ɢ<���b��)U�yB��9��Au�p� �Q9���$��H�9�L@�x�$�Z�X7_����}a���h��G2���s�e�n�������m}���-I���x$��)1�t�d�����N �& ��g�/1�|xQT�"�2���F'����c݅�jz˿��/��o/	�{�����~U��
�)]j�qo������Pa��=};Vgl�4���RR7���Ɍ?���A