XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3��EY���_���'e���t�CYK�Llf�2%LA�A(i�b����gtI<����+oDtDMۧg�fp~P�k�{w\$��k�����Jȃ�r� ɵ�@*�x��DrS��-<����y��0��5hg�õ���jMc>��T�`lѡT�:".���m�6�C��A��R�(� 0)r���a-����cs�K��n�A�?bΣ�kq@�z���2�!:����Լ����>�:�#R�1�'���V�)���U����y�T���C�D�R4e�.���U�ody%��CmZ�\C-s������Kר����&
�����Z�������Y����5h�Y}��h��l��j�}m,Xbeq9���6O�_��2p�N��:��9R:��5�#�0���}U�˗�0Z�t�������O��D�aA���7�&"���"F�OdV�����^���S�PcF�}P���\��d�`"	ذߜ����� �:�P��T��N��$���a���ܾ�#�a�����[v��p�Z��U�n /T~/(U/�����z�)�:9^|E��k�x�%}{���O	�:��좨�����[;�0�?��	�˝5�.*=�|f��Sod�������C%��{T(�3 >(�hdB�$9�_*ww�b)�	����yY]�#J	���)ؐ+�_
j�BY,T�6�եH��4��0k4N����َ�c�w֛�������[���eq��T�/}$鵘okbXlxVHYEB    1795     7b0Np�e����j���b���~ ��cj�K��7�������'�G�X�]n��p��1Fypבo`�����Y�E�X����Z;��.��=	;y�O�0P0y!mX�C��IWcHr���`Ca����<Be��PN���� ���Gȧ��얡f_��W���n�qC�d����y?���Ǯ�=��Q��WfWC����z��iH�����g�qi�����S�P)�:68�7���*�U�|�&���1-�'����i��|h{�:����-�?��f�
<�.
y}*�g��?����-P�ֹ��t&�1��(�O^k��a�����w���K�o,�����JۧX��ok��h�l�P���u��!��{5�x��<��1�P O$rȼ�r�xs�CRb�/�z4<+��0/�Y#Z���sE�/"M���;ٛ�*L�@��%�
A��<����b�Y80�e���Q���zja� CP>r��DT�<d�&[Ps&��+�	['��a |���Y��y�e&�/Z@R���fͪ������=N[�X*C<���F�}:���W�r֧떳�e��-��]�vL�cvh/�;i�7��u��j�P���h?��1��*��׾���Q�����&ʗ7��)��7��3�ܫ�&��&���!��~�C�?�f��R'D�I"ț��
���X�}������S����v�g� |���>� 
n7�����4/A�
	nX�:��^�d��S����.��-�܉L���}������Bz��y�UսǦ��a���5�G_Ј�#i 	�g.9ؕ��xd�U*O�1OE�>U���}�.�%�߸�:���X�?A2h���JL�dQf$C��>��yn��7��>�U5N�.Z�\����ri`�ԑ)�x��M��[.���I��_=�?�m�������S� �X���.9�l[���0���֠-� �w^7�rAy����ű)���E�b�p�b'Y� ��DMY-����^��[��E������g;�ep��oH)���P_���wT�kʓ���h+n�ɩwó��.V�d-�-�6�`x�e�x���]���Et���`�->W�eT����撗s��W` co�B���'�V���FS��'���㌨IY!�&OӜ˙^��Sw_H���!�⚈Sõ����>��sʭ݁U�1�B�C�Ik��#Z�v���-&��x�P� yWH�}W����ڬ��q �t [p���ߧ�rZ��:�-SM�\=�ᥰ�o���C|�?���>aT�KeD� ,
��{�qW�oMb0SY����+KI�o��g��+^ט��=��6?��
1I��>?e�9���I�f�]�'mb��h>nh!�}���
�"t(��/܍sS��Ӭ�2��ϩ�]qZ�W!��������0�����J[6h?�Y*EK���@��p�/�����g��a���Qd?�`���\�NP1E��D?�m&$���B= ��R����}lF�r6���L~���Z�_VcBv$"-�[��&���1��8�V!k���Ÿ�jX^�m~c0�D~4���u�������9�jsb)
�;,K0"\	�ő}v|�f��
��_�b��7�Z�E�X�K����?�|m�i�ͩ��'�R�ۡ�����j3f�(eIZ�T���_��Z���ml���И�/f�ǵ8${�,���w��<���]�/��>�@iKֿ��lӛ�\n��h]ա�Ucs�w	�H�<܌e��2�K�B(ɑ�WW�N��6���'g:p�ٸW�|BHw�U�Uy%|^�����ءÛ�ˎߠP�ao��&��Uq<�?v��m�.P��B�F��_���O��(s� y�RF�y�@l��$H�T�(ͷl���
��j�Z���A O�0,�-���&�^KX#��V�{c�hOJ�sA�z�\