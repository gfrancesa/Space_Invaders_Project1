XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���>���m���N�=��f8�撈m��.	p[���+�>�
 3�.���Y47���	��JY3/a<��P)� Tzw��0m�5	͐=��%�!�Y�k�MFS�~t��H�1
�/R��tZ4�ӓ����g��f92k��&�fu�������o�f~D���C9��M� �o^dc=�+�_C����v; Fz����Os��[�����k����K��{�xƳO�z)m�����C��_����2�k��EN��n	�ǌ!u� �ˮca��ݝt�);6�{z��^��	H3���|3�^�`8f�a��+x4��݌����kz��(6�G��k�U�z;JVD���3���eK��:�B���-��DV7`T�1���*��@�"�7'|6ʶ��?�k����>�2����/Œ�siuOԺn�~�ȗ4s�	U���3Ͻ;�~�Ɲ�q�;>(u��u8k���Ozz�rK�%�JWB����yK?�v؅�Sl�h�7"�O\#)�D�Ԅ���D�/5d>�x���.���t�o����)�,]�	+���46+Ρ�#I�_1���̊A5�Z� +��5�ݧ��NM권a��*���)c���-�o���k�����+nK��/�����H���&i���]{����Z��l�1<��n���^>쭬�.�8ǶN��$�ї>ƕ)�'邻WYd�U����ec1N-*��^}�CJ��-?�����I�K�{ߣ?��Ҩi6��XlxVHYEB    5e75    1150|����I���ͥs�m�j �q�2�L�Ǔ����_5������,���2}�}o�����i�R�H�jv��v������\���
<f���U���Ԏ��o��<V���O��@'wf�,���;�ۥ�{��&�6�;Ɠ�����_Y<(���P���M��3��g�Q��(2��u��a�f\ivg�J�O�w���es�����
�cFT��jTj���xŖZ�:�vvZC@¤�*�k�%n�:�g��ϩ�Fφ�����L��VķW>�}lڽ:zf���WIf�Q��E�O��hF�vG2jM�J�g�{�z��sg�%(�l�ߎ[}X�я���ȉ��c�C�Ҍ�I�X�ҿ���d��Z+��]q����g-��T�5�AOJ��~�Hi���oͨ����䋃�w�O���;��k* �yZ�J��<�Oϴ4������ڪ���^V�j��zQP�+<|��� ylI)re���@��5EU�È8'>Я�S��䕪F"DS�W2�3~/�~�������}�?����	�PQlɣ�%�S����Tl���S�z�l4e��jy��r�$`lS�)(ʠ�0T�x��USBYh�=��ޫ��ÂV�މ��^8E��K#��l�)�<%.b�mU�,�4�������p��dl��ʪ���V��Q\�����f�W��t�h.ۅ�a�]�7=A�nP�۴5\88&�dT���rz���:��9�\ԉ�����~t�����x���d��:�	ʱ����̖����oV$�K�����ap�
����4+��h���sH�M���'<(sT��d@辔�p��G�h�hg&k�H`u�5o���ؒ�J�-l��9�	{]��4��|�JۻNH?c{PcN;Y+��x���5�b��i����W)�0�:禕�G�粒f1�[`R$\H0�8tb�����,�6�d���<<�K:������ӄ��F�R�g>)�i�}�p���jpAY�wv:� �q��(Z�/+Ӣn�
y���Ϝ�HX�G`	g��E��i���(�7��$)�>]��*^�dpeX�%��Q3�̀�0��wx�7�'�4�E�d�lfVe�ժpe���w&i"jq?/$|�z�d-ۏ3�t�^�_ ��`�h�+?���g r��J~r�K���V�ц΢��.PMX�X��)���nhJ��9)�R�"��M`���mX���ע��c��-���p���u,��\�S���:嶉l1lҰ�z������<t�*��L��,t>5T1�%���Z58H˸�@'��go���B���K]�]�b��Smk���5'�D�ġ�x���G��̰@��G&�.t*�9�ľ�l���ҙv����.X���g��[�|CLľ�B�h��D7գs�+�U�y���H��F+6�)�E�h��5y��\,�����{7� mQ��X�yb�<G���2p��S�^����#���F1~2�j�Yo�C�0.��}�m��ѻϵ��q�L� ks5�y���p$�0��볜�QWDG7�w��-�T�x�*��{��SJ|�����DHO���k0MO��2��/�kC��w���rIKL&��i�\M�ja8.22�
��z�/��iG�|�R=�_��"`�0��Ux9�7m��5�Y.��ʍ
��O��fёrb�+�!T]�k�5P�F+�����dZ.BG�/��Q�*��lTf��~B��V������̘��m�!W]�VS��]�*lx�
+��	�R�T�ߋg��)L��L������I��&!���*\����I�!��3�'��*���Y����k
�y��¨r%�wj�!kR�/�ҁg�pX-��ܖݝ��E��`;\µ�NS�eDK 7��\�
I�.3g?0�]�/q՞V�/- �u2Z�����w	yF�tY��nBZ�N���D�)�p��g-��3��m\x�$9 !�_��#$F��/�)��Ne�	�Ҝ�5�,:�u�_=�O.������;[D`縉��h���4[5z�H�І���t�|����#�Q�)a����	�9�m�w���dn�C�E'�l\�̆o���O����!sҹkE��2�f@��A�y��/�w��v���|�,�sd�a-$Y�b&�����u6��<� p"������&N���)36����̨'�bP\4��3�4��P˜��SKux�?ɭ�m�"�����:��X6�������������H�*��Ŀh�֭h���N(��M[�(�%�Cn�4�T,K$�Y!04+����ΔB̥��}��C�i���JP�6�H��2�<��x�k�+"+	,2��{�*l����e������E��R�g��E	��$+\�c]RF�IZB�ȳm�I�޽Χ���t�?����ϵB��X|��9K/#����ڱ�n�?�2�_~�>�6��5,���w����C�@{�����������`.)�ׄ!A(�X��{*�OZ������i���%�i5V�j��tN��n��[���v�b��lO����K�Æ2#���~�NM�]s�<��	Fkty�F�~�6G.\�S�'j���A��0�Χ�$�9��� >�y�Qa�t~  �!W�T��gJr��<�C��\uM>����G�҇⼪��Ő��'h�?��7�S�((�-��o.ٷ ��C���h�}O�%{6� �4�Q����l�D�=�a
x�gAG�$�P�T��}�2��~-���5[b��b�._�w�	�Z}����~i�b���_�ՕiZɜ���Z-ʈ���
o��w�K�z���������:	]���֑/���EM� �W�c*��A�q=o�&�Ƞ�R����-)�Me�@���|v/*����[������W=W���Q������i��`C�����?��0��w�M�"�@�,�0�+��b`4����1�����!ƣ5$��µo��ԫ���4��V0V�W/�l�^�M��ځ�z}��OP��B`6��'<H�
�å��D�j/�΁�'��^v���]���S-іw&�v��=uoO���:j�3��${���s垲5��j	�@a���kz?'q�y>��a����r �*�rm`F z�V ��\rA��S�e�a�NM[�%��) �k���2�+�%����������s�/�m��wT��Mൕn(��&_�?�v�ѥ�|��Bk��9�	�W/`H���7DB��fa������/̘������]�"rw�-+Dm�/����{���s*ԌߎU̴&�T�d�qZ�},_�ե &J�Z���m	��"�l��1#Y��d��|�f�^�;��1�o�AS�l� ��� *m5�Ԟ#�:��i��dQ�f�_4�HP�d�q�Yeq�_g��O���W���=.���
jTrT�ȸ������Z�k�J�p��	�9g�j��s�I�s�Q�o��J����*ظ���zyNf9�������m�x�P���/K�@ %ek�K-���t�DM��P�P�yD�:bor�GT6Mn�n�}I΀)����'t��UT_������O����q�U���'���8��������E;򣊔�+�	�-d�3��[~k+]��ؽ��$dib���ك�n0<,]ɏy�x��K.��r�^L��-�r3VA/I���� �����1A&��=�k4n��`ܮ�����A1�@r����3�2*P���4��gꪸɲ�O)���F7#p�dD�Ҩ�x�O�1�.�����D�צ��
p�3�7����l��O�$�vncz��!_�4IA�o��ai%�$yZK ����M��J����e��h��pH�;1آ��A0��U��M_zA">r�{E}��f����ն^u�YE�����3�q	�	���@�v_�0G�����Ҫ��t�a,�9?~ԓi�/
�;}�$�rT�F��r���Ig�\1M���ݵ�Ʒ����u.MH�wf��#v���S;���������]�0�=�V���_㖃��vV��3���5v2������03)�����ܺ�S��J���$}>OHn_)f%�Z�a��8i�І�c�U�
B*�S����LwE�b
i����`sD��X��k5���	���1������}�����>�vx\�*�]M��lt-hB�`O�~�D�W��"oS�'��RW�ԭb	�ײ�G�|[k%Ƽ�,-㭞F����ga�[�.�� �[iB�_����͢��&�.}'G�B��7���Jy=���q��� sT��{8�c	C�}�?�}h�z|���d}��ƛ�{ۙ�㎈M�����i9�fU՝�������`A,�:7�W��3��x�v�7���t��Y��yǇR���m�