XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����zt�I�&ܐ�2m����̺��f��@��d�4�eBw&5��6�����,�d��ꉲ��M��`�P��5��~��o��0�tEs?{�p�n�	�Х��xm��*���C�_�]8;)�p��R[�a��O�0%=L�=��^�2���"0V&���R� �squ�aa�����_�<���tݞ�Ë��Թ��|H�}�h55\���Os/���7`���t߿�,.s��`�9��O���/yL�ɷ� g֮�c������>����v�!V�m�k��sQ��{#�`@)����P޹���u !��FdW�$�,|TSE��F�Gp�3��/P<����]ϒd�P�A.D�H=���H���&�ҹ�ϱs��m4�G���h*��n���c��ݦ��~p�h
��k��Xa_���զ��Ҍ��o�����q"�ڋ�FYЉ���{7}�����{i�8�����X�W�x#�P�T��w&�`�	���MZ���(>F�t�@�ί5�$d 0�,�C��h!3�4��m*�ߴ�����JD^�h{����0��~�V�?}>��O�}���(���q��Wݰ�^�SBy��Gє$������W{ŏ�Vח�\1N��{��	�������MC�5l��?�'� \ruSme,���Ƃ��Z̠jqw��!��S3t	v�R���f�E���g;�Ȼ��>���Me�eU��w���P�.w{�s�r �)���b�׮мve\3i[�e�F�źц|XlxVHYEB    6e28    1620�T&�U@<��x��l0':���H��B����-�\�-p���!"���b?pad�z�0H���PĶ�>GOFAQj�y�3[�[�������gd�`x3j�l�s��.�J$����� D��ؚ!,่�+ɋ!�ej���p��4v�����-S���(&f�0V*C�C+�Ǡ�)`Nl�xe��Ơ�5�}J�С_�k(Z�y��ȇ1dCv+Z���O0�ڰ�4O�Ljm��{�F}�n��#c�����6l���ӣu���*��\UXy���M�p�����j?E�H�(�����HV���=�����|qъ���F��&��u� _Ɵ������u�,�}6p\��+���,��h��'��k�PǮlc⢤��M) �d��q�N��>��.��Yw�(�8|-{^����;�����2��@��[<J�d����X��En�-et���A�(����nK7G�-�/�Oڇ*��}��6:}���g��g��k;�ʌ�R_Xh޲T��\�	��^F!��ͣ�>��W�!/�(��x���ũ�YcnN~�YjgYN��yn��,� ����o��2�.(V�Hy�Л�/s�YVg�ئk�!0ZC�q:��a��aG��xTz�R,�`���`�;A�����tnZ�`p-w\7X�a�`�pӍS��TN��Lt�����
�~�����1�9�wɘt�*��<&
j\�d�J�`�âށ�/���06��Dh�h��v/�~BѠ�_�A�+̔l����m�I\v�T�E݃8����<�L�������?aU���QI���ˎ���7uܒ�ǈ���ggH���,�v�"ã(_��7������M��B�GR�&
�x 9`V
����gPU��<'�?m���x����}�U��V�)3G�n,�e/V��ӀI��dZ�?��_:�����/�d�]�=X��6��C�b��Tsm±6*HSf*J��Y
����g�P4S1�/��7�8���U$�Sj-T��r�㳭*��J�B��
tz���`����de���h�\#،��g�l�P8o�����1D��g��_��ǹ(�E��tJ�m�t5�<{t�:�����%LqOC_��rjb���toELۖt���)��kn�Շ
݃���j�0K�@ϒ��O	j�
�T`#���.�~JP;^"�%V,¼n�@�8����LJn0��l�\�.G�Me&�Q.�гT2^�%A���I1�A>�:�*�0B�	_�d���g��B<(�U7�6�2"�:�Pxc�R���GԴ�X�ٶ�-7��v��\^Q84�����fx�)�T7p���y�T@�i�S@�L����<�	�
_��zd�:N�Q�KE	����oRʶ����R���Mi-a&P�ND$��**�(��
�<�x��P�B��qN�^7�h�ޥ����v
soLUG�yܬ`0�wp���GH�qzB�����F:l$f���Cޯ&2���M����C��m5!�b���S[�F�e��\���~�29K�Z�_O"]�c�����������pi}"��V��~+���m�ݡ��0
�ҪF!4;�S�&Y�k�#����o������32�f������;WK\�EH�н�yZf��&�2��T���0=�D�r$�"n~��G+���6Lb
��r������lק_�HԺs�p�X� trI+������y�aA�G�706S�Ɇ�^�.�Q'�����1D���.(i5U���2�Y��k�S��8d򚬞ޜ���Ι����è?�;I�X���(��ܯ���Y��a����Z��i36f"�Δ��Vu�A���#6oڙ*Y�8Q!�Fӑ��xf�s��K�1���t�ٲ�f�u��.�u�	��ݯ�� Q�����(A�r`��,�=���OPa��r������n"(�;v���d�b��$�S���&<��~ҏ�E�˯�됬N�����^��)�� ���B��<�虽�������b���@��
�9����z�KG�]-��5�/*%�V�pj=��!�΂\˛�Jy�)iV�͸��嬨�1r�/[�f�.~�����A4�@�XL����΢��V��&b���?E>�H��t��2ˬ��/51�U#<R�����1�1�Mp$ml�o/�%�3��8�=c�8R0"�{�O����B�yA[���K���
�lO�:�
4޿�QBD��_k�����Jr oy���K� )���u��'gt�͐�N��$�뎓2��N3U����~�}-װ�I"(0J��v�*���MUK���ٺ��K2*��Y�Ջ����{c�˷�����M���IЮ�U�2rzXeW�]z*C���iP_��Y�N�	g�*b\��l����ݖy���˭r� �F�/�L��W�}90DYg5����ZU�����P�e�f�\�/�?�S�@� s�>z��hp]��D\OM��܇L X���W�W�XT��ա�ǰ��_:���tG�22�g�h�9 ���"a��<��&���6>����������\�o�����Q������s���m�Pl�6���^nA���홅�K�$v9�+}|���G
-�I�e@�{&�o(SZ���.��C��i�|a�x"VIdL�M�҂�a�x��$�Q3�ƛ̊�8l��U��$�\x	��s"7wem"��9R5ْx2�e��>'��"��'4; )V%xJ��h��X��/�;2MX�Ap�����Gg���[h�m���j��6� 9����*��
�F�u3�.0A��7abr�	�=�_�#M%���w6K�ͮ����0���j�^kq��;0�]���F�`��+g�E2S�<q�w��O����� �s=� ��'���m�C��+/�,��V ��N�k_�K����#|Q���կX�d�y4�?z�dn������r�]�iC,��'6���%�6�jH��@��;�\C���:�b ��ف����G�aOԜ?'&Ƨ{����<�l�Aqױ��W#Ɋu�+k��tf� lS���	�[#�&'�>1)�
$�c5yx��qOe�G�Ps�`�䯗�#�a���Uк�jxi�s��HD��꽾�Rs�Gx����K�9�[c��}�/V����߆��$�JN.�R�Rv��Z���AB� V\19�sJ�D&.Q8ee�(�[��Ty"� �9�m�$�¿�˵�����&K���*�`,&�<@P&���h���UO�wG��V!=�j���zNS������L��3:�ϫlRop\�_p�k�B�TU�r7vJ�@��:�7l6�͐4Q1�F�X�g��Hl��Z=� n�X�����!��X(@_�X}�s��cd2ԓ����pP#�-[A�ǟ:��;14B��� /����e�7�Ւq��#���h5�����-��X�8�^�+g�B���{��;[���m�1�����1�'ˋǧ��=���<��j��*�XX4�F�l��������z>��Q���~˲�_0��\;�ƧSAՉ'���D$����r�=?��ϛx�JZn6i�gB	`f��u ���nN�fϭ� א{k���
�g'�2�_t>8e�z֟��/�W����-���8�;�FLo�Xf�QD��H�ֵIĹ�l��@Yl�}���A� �_�_kG��3�G�|�U�T�}X�E����9�`kˊ�T� )�i\C���+�Uuz�V��D��3�#��M$�hO�k鏚��ԧzOm�7�M2k��K̇J�E9�M+��_�QJ!�&q�
Oҥ�4���z��O�c�o���_0�Uvk�!�1�-1uB�is4f�zb\��Hs�/�8��n#2m^�S׵�^*.�)��;��޺~>�Z�t��A�|�p��G3vW�4�'Ⱦ��8&��¼��]�2��R�u	��� X�5��ߕ3�`����m^�N������>�C*��N�P���'E�f��دOc��z��*z����6���;���E��
~���3Q2��)�~�MuW�_	��G��y��xUN��0�R���*U7 �F��U�1�,Ȧ��W8�o�GW�W��Y/��2�n6r�`�+WԷ�1 l@B��L�.�����cC7�����,�~��|���Wvg�i'�ۅ9!��(V$#����v�ݖ�eb�����#ۓ���!$��8J��3Ǥt{3��نlɊ�R�~����C"��ſ�Ħo@׀B��50����n�O6ڏqz�l@jV����(���_�z�#����RoJ�}�ޣ��i�=��#��Πb#���*z���G�6}�k8�C�d�*0,m���8.Ϸ�/���*�(mކ�5{�'�DH ܒ�\V�����z��1C8�:�0 ��3��Z��z'��=�q�E3� O�]�U��D~#ԇ#�����R;��~�V1����!��~zz4���Z�z�+��J��Sش�D��/օ��y�)w���.~}P �2�ۻ��W`���#í���L�2�\���O/�a�ސ��R�ɤ)mC�c�RG+j��7��I�|���o��%�4�g�h\i W r1q=��(��ǧ����:	[2��ta�����]��T�M���̣����XxQV'M��a��2[��5IN}3�^�����n�ܞ�k�A���\����� =n�Z]�"���㠝 ��8��y�F`�7=n�}I?��<�3�_��䁺vŘ�'QI�?α)iȆ8&k��ӣ`k����@CR�}���2
����=0#5��x��&�N��Q/,��${H�l�%��d����<��>T!��AZ�R�kwPN�p}7f�� D�H�ǆ#Xe籐��:��>|�;k�yg>Vu�	;�7�ɍf���(`v�=�ː�Xv?'�	83CӭJ����Ѐ��5J�@|�L�}6X]�oU��rw�o2��=�ew����u�:S.��~;<,Y)�k
#��˜U�.g�� w�����)fr�&�.�i��_pB��t�7۬W��IE���q��S�!����W)�\E1p������}���_�|�@��� g+l��~��۞nB��F�4M�5J��caj�WC^O�N[�==�A�鴟�qFMU�0xnc���ᶞ�3)��CVޔ�c�F�����*A���H&�tq�h8X[���#*:���^�2��#��ZT�:2k~�U��$����Y��G�u��㢺 ��o\��6+�����6�n��g<�5y,�y�.tp����f��d�ԫu3��<�U��7\2��X]�]`��&��/����N��,�C����Wwٙ�Ie����/�a�|t1�qY� <~$~%�Ԡq%;)��	�7p&���@���qWIO���I��}'�O�(�����N+OHrO����z��P
zϑ��h���_9��h����.,�5kh@h�f�L�՗�a)�B�e�QJ/�d�JU�/�����Y����
���X�e�C(૳�0�H1�o��-̵ۓ���{/Q;I���3$�ZA��׮�
hW��)�qՙ� ծ�R�:���˭�������Q��