XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[�ct��˄�@c穳�{Rg�>2��� ����� �2=��Y��jO���þ��x���$)t����.`� �A9���Ϝ-�W_�>��ՠ$�Th�MQ���"hq�4�ja�㒆�݇@wZ>�'�٩c�&���O��?�� ��@W��c���(�^�t�9�[�߂�/R�eUJ���>e�O	��H>U��00�6����d�wx�F����M���A�څ���f�Sh���������\��m�Yk7H\�Td. ��?K��t�p����3���n�,��ξJ20�
��o�3w0bBu�1�h�h��:`�sN��+�� F~�FĊՉxN�R/aZd)+@��<V�Mi�LC�7/B�坚G��U�u��T�-�����ٙ������Cwu#l��� vQ�#K�pKCR�A�d���3n�Kepo��0@^*_���ч���Q[X
}�C�����sۡ��R��c���5���_T덷�3�šk�6�&���-RB\�Ge
@8��kQ��o�&�A�����k�$w�-�v�@Ҫ.��k6����^��o.G̬��F�ܕ��G����dŠ�>�HS���8���/����-\3 ��yP�_����i���9uA<��V�X�S7���C�u��S�t���\��SD}Z8��̡F{���jf�/��r���Q�Գ�[�'�O4*� .Ya5�
���me�޷�jxh�"�6@���N�Z��dY�G�XlxVHYEB    2bba     bb06��"5L������:�a	4SQ�B�r�*�N��/�s"����8�z4ϑ_���)��I��_q�e�Sh���O�ˀj�������3�K	�2��y�*�&��������}��ָ�?0���ZZF�~�~鋉�f��uA�0qC� W���/S�w�0���X�"4��!��'����k�A-�q�G�U�u�����J��G�4��tm�CMQ����W�ʘ�t���#z��#���+P��u_�	ݧ����#?(���l��&�>]��t�4J�Mv�8�%��md4E����uz4]��PJ�oÇU�ZX�H[)��C��g�u]����Yc	���������\�e/���9f��+���GEv$�1���KZ�q�<��o�ϐ�)��A�H͇�l�&X3��\�iR�\�\݋�����ҌГ̸.�R�㬿�T"2�"���q^�����K��dq�2���՛�8�\&ڙ�S�{qH�XV#�iN%|v�1�0�Jr�z������;G�\��rZ���E�T7���q!��([;�b�U495H�jD�@�m�$S�\?�v4�����Tе�Ⳡqu�'-H��FU��j>�iݹ�D�#��ED����Mq���������^XC�#� 8�1�![��1����h+#b�:���Q)nr>��ߎ��$>�B������^��鰰9˯�,�t��֊ДN����7���}�G;(�?��+ƅ��܍�J�g��$ru���*}�$�������/���~B�3+��]�d�k\)�h��w� ��Liz|M�����;e���C�;��	!+1���=�Ϝ$9��x�}l{��5��QN̩����U
�;���c�I�:�ٜ�8�ͪ=�4U����v����9�h*h�s�*[��5��i��D�������c!Z�=���h)��	Y.s�ԍ٤v� ��l؀�N��'?�e�<4΀� ����6���ο��u�s��5>�W�e^F=����F���F���ʇ9�N�J�1�%c��"�obIJ|E��ZPݼ���
������"	��a� �d'�%_�^��'��uCh��u�Nm�D� ���,K!]Z9Rle��@A�	�4w��]�"���\�����va���Ⱦ�(Uشа�<���G��W�*Y񬶴�ó���O��]������]��`��o�-�k��qAa�S�D�5�O���|���/�):lC�����
�nHf�<µ�tFw���;]�˩�yM�B�X�A�Lװ���1r��~���BKO���.�d�v���f��NC�=��_����FAR���ş������+�V���2�<���[�$�#��'#&�������������*����I"žB�v�A�Nͥ�W{lum���(���M�GP����'�Ǔ��A�`=Y0RL��-��o�Bhw�����2lX�8+R�9��L��fCau�z�ڪA!�4{�������nn&O�̈́��"c�Ӥpr��!S��q87�d�#9&�^=�j��.�I��� V� ���STUG֗<���q��p6{�[���ƭ�⠲J[nGl�"���{�U��^��5E��o� #.@0��4h�k�:��)�Z�b%槶J�h��}��H=�%D��5��F÷�B�����_t�����W$�w<Ҭ�@T���"���:���DG@Ȉ�������@C�j�8�=��h-4N��{���<��g�ԺSO�<Q4���c�3����������׳���O�E�I�ʗ��R�i<bvZ�]Ђ�_-�Z�	W
5"�.`��,t��
8��Y�=�#d��d
(��x�3�`�=H|��m�n鬥e�&��e<{�窎� �f
��w��P����5�u�Ń��|�[%�]�6GVof<�sf��1��>��{g����Ў�H���p�ӄ����DV �\N�<z���KY�0S�A�4x�/��&�Tc�fw�:V��r�w��!�#`06����Z�RMqV����3p�p��a!|L�U)�[g���.楨�!�<�Qh(N\�|�ֱIAA��,f	�3��<Y���.�#|��Ӊa�B6�8��%�$aдP�B�eUf6�d��ib�{�ۅq�<�سAwu���%G�k�_~嘎����Ðgb��!w��ww��������ԗ�����y�cU�!�(�����	�x�%^S=�J�$r�C��Lp�f���*��n��2fx�F�0�^F] ��C$��=��G�y��z�� �%��\8s�j�W5^���7��)̊NK�$�F� S'I�J��K��;�*f.!��(��.i9�r:�
�����DH��#��z'���K�JB?��p����i���g�q�;��ւ; Gw����8ٖIn¾f�	�He�g��9����>ޗ��y��pIZ[hv��MHB�[��y��������c-�Z�¿9�3O@���8�E�^��kXE+��Q�ȼX+ۍ89H���8���w߬�ՍJ:�p��i���fz�DR�'85g�T@M�廏�p��*�K�ͥ�_V��xH1��0O¿�e�9f�7#~q���_9b	��5�v����{rrq�8&%�x""#z�������O�̨���F
�\SH%�:�Kd����t��r���.ƺm��'�#�X���m�#ei�oBL��#��H��~���_��K?�����@_�eP���h�H�~B�`��Bu����V�����6�4|,���<+��	����>�����!���PA9�ϟvZ�P�S$�����o�����0	|��9�Ȅ�F�)������-�wɺ�j���[1��*9�;�R?�/����vSW���#��o�{�~ƪ!��pI{��_l	<BR����z�PN�dy����3����a�@��]gȻ�X�B����