XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��j�re]P������"��ID�q,�d�!�^'gp�����Z�p�r�����|ȳ���#���+a�������2�T��c��/��"�)�w�9D�*��J�d2�������ޣ/�O�����η��!�?O��o�[ڑi9��Sϕ��2�_��^�-������o��}��ؘ�G��m�~#;�覵��-�tj��+ͨ؁
R��C�
^l�nG&�޵�Sl>Y��W�ͻ��%�&�S�^�سr����VA����zd��F,��:�S܀�`�|
�)����(]E\��G��V�E^�ɔQ��z�y	�J��!ݓ=	BAjh~���3�I0D�%"f���;GЕ�2�ғ�"Yn����ЙJ�|v)����lY�u�xY��ˡ1kZ�}P)��R"@	RƫKԺ���kG�����i͌���#�0s"���'��s�C؉Ctj_�A-7��~�m�K�ʴ'�bL=�̄���$4Z@�YQT��H�f��H�[�U�N��'6g)��]�u+��X��|8`@���Zg�i*u��ukY���%���^)4[�qbֵ�jm����_�4~-�m1ɂ�3���0[�$2,���}��q|w�����J���z�v����4_�tp��]������������S-6�E�n��|a�� `%g1�C�N�lc#��Ȑ��NB�
���6���K���C]���0��M����kY�&�!�uE]�LR˖C�@fŝ\�DV�f��XlxVHYEB    4ba0    1230������b��#T�e�rtN��t���f[���wn���߇�*�#�ςY;�q7�8��Zd��=����
a�]�����b.����X)�>��I��:Ȯ�9�O��B?L����%5��I�Si_�	�̇|��c��q7���ZTx��xE��ϋ+���J�>��Xb�a�w��ACI&-�C<��IU��3q։T�����eq���N\i}�+�p��r���p)�O`��1���]nx���&�Bײ$�B�����y���xHC�VP��@i�1�/��+#��K������]U-ZM^"���A�����e�0�H��c�I��x0�����-�B�A7��Kj{h
5�Ȏ�-
 �a���S��_0v�U߶���
�#��v=�r�ʞ�%���-V/.sʣ)�0�\\�*��]����="�����,a�փ1��#�Eᘒ�N)_g�6�N�Z�����y�uS��tC�,6��V�k���]s��[�Z�_�u���9�&U�Ӊ�i�N��v���(�K�`�-vY�P��G\�(ogִq>���cw6'2E������F�qzt�<�oM��'��:���j��vξ�����=)��D�LP(El��?��Y��i��c)կ`�_�挢;�tLc���Qt�{V��/ψ�*�o�Q�cڢq���񫬁cn�����v��\����m� 8%�j��îk�_hM�t^�u9��kﺐ���#ѕ���� ־H+�������7�&��c�'2��T!G�MB˟s�8U'1�?ƥ��w�T�c1�X!jA�w�4���O.��A^u��d���z�i�{1��HQ��槢�8���I�G�+�$����Y%33��)D�?e��vKA^Ұ-��f��bb������s�����D����m�� �;�`����T�z��T�E�S�
7�	�O�f���j�;��$\^c<>Z�[S���jP_MO���"߭��=<6{��"�1�s�j���X838�!�����1������:w'��q����`�^����7���XJ�� ��b�P�����c������hz�+�t�1i��hFR\�@zF%�H��#��\�!`�J�rc;�5k�-�j�^K\w_Ax����Sg�5_C�[c�o7߁��b�C�k��ƂrK,f@%+:dt�3*���Ѡ��Jw����ʃL�ش�P��>T&�"�����D�ԫVl�ְ��1�y�#��0k�</��g�6�/"����'H!C���
m�&�g=Qg%wyTNA"T����@;���L>��=Y�q>����]�t|{��0�TK�2��Ъ��, -X�<mA�U�n!_�M��7�L���P���4����8mњ�Ͼ�^�@U��A����y�v��G+��͋Ti/q�~Α�z{�S o�+[u��[n�G�-��T2�؟�ÔZr,��lNp�-���v��8�I��lFPNhʸ�k4!ʞ����t}o5I�9;U����m��~�����Ŵ�Rc���c�e�"��A�Wj_��@w�Y+���<���/�z��&[,�G��n�L���M�K7��	N�:��m��g悄��(��7����ޖ��� ��;�Ts�TE������v��zx]���΂:���\g�f�T��b�_˕�!)�((�t�M�Cuյ%�i��^������@���#hە����������S��&&����,bTlH��E�+�u�Y?��u��O_A�B�5�<.���/q�V�t;�(D�ttT�މ�l>�q-��;��ɧ��m]9�Uҋ�F�uQ=n�y!3���RRLR%��v�U{`���B�]�;�^[�p޿^�ڪ/�J�IV��ցSy'w5_���KH @�[���w�8�n�3�b�a�eXJ3J27Z��Q�*}���ŋL�B����4;/y�&�`���P�Dn��U����q��x�n>^�Z"�X�C��tĂ$����8Dv_OrWG��RV���n��)�S�0fɴ�:%-�|Z6q�&s����.�r�{!�t.���uݬ��9�N�  ����CzPS�7� �I½�5�8!N8�/'`vC)EN\��e\w�_K�@�j�}v!nўV,�}�Y;8@��V�f 	=X7�+�x@���d�I��^àq�P�B�\Do�&�9����[��:*)y1��%o1�<73��d^(���u�슕�	$��kZ��������*�-"�-�'���Ғ���n�8�f��+.�&���Uԥ�����>�ʋ���<�������Y�����t��g�h1����W�}\�5yn��׉� �Q8�x��ڸ~���@��x{�\�`�V�_(o��Levt��9���ɫ(O�>��6�H�0C�u�"�����(�a�d8������Cܺ�%�g�6
�$J�jT_TZ"��a%q�\�A��#`D��q��۬*�ޒ9�#��ԫվ BAEr=�S.��A���w�����Ǻ%v���hә�Ai�JO���=��2#ѠCh2���gm�rS���˖(��t!�*썏P��Bq�1/�0��|b� ��[��{��� �+������¢�W�Jk�T=G�$$Ntr�@d����t���*]|#0��,gg0S]�b����.U�����ߨ,�9\��C��*��sE��H�V�h=AIw)�JX�|kn�T��}	 =��a��f�]�X��;V�w� o{�]�کRF P�D'OǞ�n��/�r�ke䎡Ǆ�rl'�b�|G`��	t�N+��VQ�"3��|�9O`Hy�����G�Y�e`i���`b��ՒFqu~�Y���rB�^o�$���h���Q�R����m�EՅ���)�w7#E�<���,[�^m�7R�,D1}�i��,������ y*�!Av��AJim�_�'��
sKA�����]¦�n�l��d�/?�z��f@���H�H�g%dF�*5�h6$�kU�7��xl�/��Pv�c�*X"�vK�b�~����֥�� ru7=Z���*��5G�������-�C�*���q�.�����:����l$n��<f����=��߉��R3�.���@&���G�0�����n`2̾���29�VFE8�$��!�1��'�S/�b�AOFJC����B�di�qQC�3gv������^J-N�~��&�?�����.)�ڡ�E͊/֜��#��({����Q���Ú
߉�aL�ԻO66�{�@�%��0��2Њ�D"NT�om��Y7�? ���`ԔJ����xDw��@�ml��|�zs��r�-/M�^$�9�
@l� �KQ�U���pѿc�"����
�(�;a��쫁�&����E��pY����Wht��l�������hC�_��(�!���y_ʨ���� ��eӷ�S��>lr�'D����r��������6�7��_յ[(a���4hiNQ��"L�أ��Iok�8\�4����˧^�tzC	u' $F5V�7[�l^SCEi�_o��D�O���Pܴ��07��;��:�<
���h�
"�ɝ� i�����#�e�r�E2�F�Z��14f#$�0K��Ư7x�)ÃA�
����8��Zû������f���k�~��?+[��7]�U��0���Tg3�H���ԉ�{ɔC?ۅ�`���!*a��ST!����T�I�}�-��Ĝ�Hk�`sQ�QVn��c�ױ�d'�7��2z&�W	��ⳝ�Υ��GI�T�H�y;4Zĭ��[MP9NQ���e��F�OT�g�{R\!�;V���A�m��^"
��=�s�Q#-�QԱ��R����i�P�<C��4�"�G��`�0o��͟Z�6,��������s<���t��`A 8f@�����w٥����s�������IE��b��sPCJ���_�&�� r�0�_˕��!���iXO���xj���»���<��gW|�Cp`�n�׊iU2�+,دܮ�/�W�� �o�L�օ><��h��8�r�>�_*��. ��&_�_7]��7��������W�+�X���+f AK�����^��h}6�Ql���k��= =��+
bH��MC�#�U��wj��R�pO��Yڂ>j횊�}�%�)�;�O��l� ���*�ѳ<��W-��2���n�,�{�y��k-���m^�C]�q�u.���d�q�BL�k(Sу�(��\�ޛj��VT����L�����i�+AC�F�Úe��CzUFx�&�c� �[�iЭ���x�DkAg���� ��8@�kG�a��� q��܃/�s/|	f_�o�#g"8-�[pɇ�߭fwAi�3�TC�z8*�0�]�HX�����9����U��� ��x~�t�ĂW�!���X�УCH*�k��3X�*Qx���jb�s��t��y*�>D���@���d���ǭ���L4KQr��X�:bZ����neV������z��^*:��aX�#*�B���'kpe0�?��<`8J���7&v��5��j�������+�M +,J���[�$�2xىaݐ��q��=s��;��A�hP��ռۯ�� H4؄�Ei�J��yw�GR�