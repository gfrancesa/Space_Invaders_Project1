XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��|�|�Ư��L�W
Ň�D�Qq�Gώ'f\��k��T�ȭ�m��¹�1%nWM��Y������i:s�|�|�уg-�7��G0fm�>R9\9�3�}!r����y
���a��'C�'��:+�{$�ݨM���q$��M1Ok������[]N���c�0�ݮ�ݸ���|\/D��rt:��{�W�=��i���f��W��Q:�EB
9��ۉ`3/;y�O�B�R�2EEpx��MB�6E�׽-�J��&��r~\�ԢΩr?��τ�소����P���`UL�0i$3�w��t�֞�w�0����;���-�)���{���Z�;��{��*����_K>^�Ii���e�A'��p�ˆ��|l�^C;0G�˭�_8\������".�yfQ�����8��'����d�fVwf9LAL�����g�M7%S��N��/F���0ʑa��H,���G����y�ޤ16V3�L��o<DY�j瞪�%����h!Jn���-�r������ս�d����H�W��*�1*[��ݲ���
g���8�P)���i�Uj���n�)�\r]{�~Ǟ��ϲ�������<Ľ}8��mΰ�a@��D��r�bm���R�ka��?��W��� ��tzϚb��O����,�%o�'��\��t;��4&��`pu��]N)���)���	>�i�}���*O���l�*T��1	꼝LŻ��/1�T>C�%n��N�mx��s7�V(4|��a�슈 ��y��DDr��XlxVHYEB    4013    1050���/حu$�5a�h���̘,���$��&�s�\+��`�DM�G�a�Ɇ6Q6U�,���f�ǑN.H�jE���_ߡ5&�t��@�3�֛�J�ծM�䉐c]	�W�V�`D��?��z=�]
�n�O#�[���f�eX��d�}��e�&ť�Hk��cѕ��I���q�V�*�9Y6H>�0�:�(@"M�7�F���,���]�Y,WVL95/4�~��(��Z;�����*do����x��z��%�"��1��0�MLOv��h(�@QCa} f�����>�� ��f�;�ڙ^]�/�������ؿ�<����.����p�Z��d�$�Rl�g����O�:��"�8�~�N!^Γ����=m[h<�n�aI:Gِ�CV�̯g�V�"��׬�:��v6`o嗳Z��cD�e�z�w������<]A���.>'��Vq;.?��FF�۱��w�-��E�w)W�gE3��|ׂ�M�n�`~B����?�VT� 2AiEc��]�!�kXg�?H�"7��L^��+�y�mB)��`\H֝Ol��w��v�2�c 霑�T������&���	�Z�����;e��55`i�<�� �t!�{]�*�1��z^���.n�@AŏGE��kY��+�|	���+�?v��k#g�� ��&S�;<_�Ps��}S��_��)��G?�V�-�2aj���:Q�L��O+���Y�����b4� %�Q�|�)��O�
[���L	1�	���,��T��	���D�Q�bhȩ0'�z'Ì�U~fFs|��	^� 1b��<?�'����:�il5||�~<�U��yRT�?�ml84��o3հ[��z{�#�����Jޠ���h|���a��g �n���q50�NKZQy7�Fb����u�Lq�i��Ş𼣿|�V5s� ��r��!��)�9Uب/�>��P}�|8*�&��2��gT��W	<,2���N�U8���P?QN<�+�}9ᫀ�
�eϷ�I�ᗪ0�>�K=P�E��3���#fZyrBSH�=��G��Ɗ���T.<A`�}��5֜�3�o7�H�7Re�}Z��o�<Ɯ'�W,Fi��)
R{�B�0���rR]ļ��ϖ�l�a^N��l�:��q���Oڊ��qCW��FP�����gME5`7��mj�������	W:K$_�E��$�,V�E�b�}�|���ܶ�~V#����!m����Rۺ>��Z���^M�w�3B3ꭾ?+��"�H<W�%F�E�P�4j��*�3�׹�4t`q�m?b
�����P¼K��	~>/M��0Bd�hbq�#}�~��/���Z��S���pEo$�����wxd�!O�Ȗ�����i�����e>?Wͦ����;�>Z����	�$��f�%�%�D��_�eA���ј!DNq�گ�3�~{O�Fl�L�c!�U0�l�bJ�EI���O+�/����t7�8�AA(�S�����>=�l��s�,�jB������৵�0�'��>�I8����Z���B�x�'�IF�Ľ�Ν���t'�� �6e#�{���WN��&#W]'c<?B��G��r��8�&��ش��P��!q�^�ˑ݅�*�B�Q��q�:^�[����0J�9ڢx18(�A�QB(�e"��vSHB��sc�W����( �����a�������0�lS�{
®.RѢk&�V5��+�Q�Ȩ�a�ә���r��c�=U$�)�����Xo���ܦ�������&C��D��\
	C��[xzI⧀l֒Y2������.���PoQ���,\5~�(�����9a>�/�J	������OL�g;�P5CNq�u,[2��g�Q�Ol�,��5zJdx�#^�S��cXw���_�ph4�s�.��nœ`�������yDupmq�c3f3^Lon�0�k��e��{SǁsQ�Dyp��������q���z�����;�G��5"~Y���*�"�u /�x��Տh�v�_0Fum��ܙ,"G$�Z�9����*'�y�Fj��YƦ �W�;Y�*����%g܆�%�X�A�C�����]��S$
�G#?B��m�+���=Y�D:��8� ��8zc�F���8tt׭Q�N�N	@s�V������&/`��tĕz��W�,�:���QH%%�,e���<x)g�Բ�%�ͨ���m;�I&~d�!���xf�Ǹ�CT�lˠwNc��M���Ɓ�$����3���;�٩�}�:9s#<�Q���7��Qk�F��Ӽٷ�7�6���fc�jf��A��
�p2)?[sB<pŘ0N�:��Gp�V38����W��/�ʑ�"��Z�m1�� nbTÇ'�5<#���fj��Z�tx��%��ױ?M�Ԟ/�\&���+��/e#����k6�o
��u�x�-#�"D�����)���)��/��w�c���o����Q(��\pߝ=�+��dI昊e��=����@r�f�s�CI�i&�K�Of�5~�A�"ZP9��=�` 3���o
'}<+�d׶�
�6��#��1�7�D̈́@o�|�U��rF�	V���Ke�*U\`�A!Z��ZID��+�薢Vӌ�w��K|�:���*!4�`��A�^+S�=)�����}j���q�*��&냙�3�:�貜7��{t2��,�"܋�JK��J�x�[�y��5�d�{�vk^��/V���)e�@8��h�lj-������gݑ�0��UJ��q�S^X��0�1�E��k�(�)l��o}T��2��k R�U���h�|v��køR���cW�����m�@����\�g�(	�e�t昺Cں��)ϴT�n��{'tuۋE���m����u��YAZ`�$,l��Y�BoH��&`�ʯ�/p��P\&#�1&���5�f�$'l��Z�� .idAJ�l��MN1���l
�6#�%B���2����x&���J�a_�I+�
clڲn~?���S��1���Uo��9w����X�{ˣ�O�Î�Z�*`��N��D��mM<l�4�P��	��1�s�Ҽh�H[[:�j�(S0��{��s����D5�6ŷ����<v�-afҀ=�vۂz^Ś���H��N�Q
Q�x�c�xG��lt8ӆ3��(�@ЁE��Y �0�~�9F�L�(n�)x�q:���n1�u�C�l��|�	u�C�(v_BPK��Wl3�g)��SMc��(̖��u���,$��L���d�Os�ɡ�R��rӴg���T	4��n�{��~ 1S;�#dÇ^��&L���c�ɒ�2`(�,�ಛ��`衧��E����x���om(��Dy�A�/%4�ŝ��N�*v �F�ʹ%?��:��'�Y0^G���L�3���CTI\H�>���e@���}b�]�g�Ҏm�W*y�u|��!��H�+����Bq#���v�3�����'u��>�ѣ�/��u<0��(~J}����=�!�����T�����V�A���P[].�ߙQ-���LI�*nE3��=��6��#s���j�"�.Y<��ޖثH�,�����5V8-Q�7%���4���Ο��z7�4�f�8���t�Ƽ�2���}N�Ʌ�O���e1T�f�ٍ�T�ou�֏fi�z�;�޽6	��&@�d�J>Z؝q£dy���"wm��f�
��F���)��[((	����jDuMٞQ]�pg�0Կ�Ի@\O;�K����h�H5���x��רd�w���j�dL�����.��V��1tN�D�ҽ�	5��k���l/y�#V����=p��-M�qy��M�ǆf�t��`���W��N���~	ʗ��}�2�P"�'�lEᐘR.P�Y���W]z�{�^���og���v�ce��󥉶qb��>�V���֏`��Qw�bB�L�����9�|�e�ͥ+銹�H��I;��u��m٬m�$S��������y��MsS-�t�VtkL�[.�j�Mo�#�D�/�e;X�q��0��Z�9�6�J�Kl�=׏�$�)i�X5�\�ɨ�a���F�ތ9l͙C��T��S\�3-*|XG��O� ��f���%yE�H���I뤧�'�n