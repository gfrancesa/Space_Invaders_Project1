XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��׈��af�p}e�jX��ί=8J���;w �eFa�x ��Ҳz��� �9��4n��HN@�`�J��椰$.�|�9e����0��lQ]]s
�������b�t�;�j���W��x��v�[�Pu�����
o����ȱ.�����I�9�o�R�I�"�qF�L5!��I�%1M	�}�U\y�u�z/����/�kˁ�~�J3���ug��㘋F�ڞR�E�n(X"�2�3I��b<���[��n*|ΒC�8�o��;������zr�4�)0����YUM�Fci�d�����$�����I�K�N�0\�w:�E�PP��.�>�bL1l5f�O\AAD�5"�J8H��f�Ln�3�ʞjS�[�J%�W.��r6��W� <E(�W����pa�]^�f\�˅9�Kǲď>������Pt���F-�)U,�l���L�"��j^�0�N>js[(䑔��<��$c+�}�>x�ԡbeF�U5���{L�b{&LJ?�z\j���~�͇JS;C�R���a%�I�o�f���]<��!$�$�_�K�2ԏu����5��[���Lm�<{�U����L谵:�Q?a'�Ms*#���M�r�O�YB�9���Z��*��n:P+_5�0���6�m؄�)��6�H#�<�m׬�xX��Y����Y�S�;�w�X�8�q^/z��V�%V͞[������ e1��+�PS�D�������]���#̄�pV��1ʳ��f���_�Oc�*yXlxVHYEB    3d5b    11c0��^?�|�C&LX	�+�c��b��]gZ�h�A�Q�LX/S��@���]�_�-5��I~~{=�S�eo��\|�!z���+R����걶̝A�b� ˟~�~�ು�r��#j�J�<��rE_����������흨�&����CQ0I�xK�����L�'����J�;����k2�j����W�ZFIW߅���X@�-��G�:�@q���of��O��iI_�gY[ʘi�'!8����]��HoP���@b�H�/v�o�5�dvW�7�Y92�n��.!3JV�z�:���c�z�U��iq)
!{1'�.m@J�]o&U&�-}��XHnf�F�a�1	��K��h$�������]8fH݌�я�#�,��HB\B���.�#��b��ܱ��6^{�֚�m/VW2p��)KP��J��@��/��~�W�!|�dL�78^QΤ�2�b�Y���������hLc�9H\7�}e��W'��ujɰ<���ӻ�7��ԋvHΒز8b�ν��K�AϘ$A$�C6�V�&�kEeWN!�$�Oxx��#�:GF^�;���vL,O|�Ac�Ճ����}Б���1"|C�"�5$I�1�մ���t��B�0�^���l��F����z@� �hR��0 Enqpǣs���z���Ϙ pf���̊uˮ�M��$�C��w���{�Ml���H���!Tt��R+��k���U=���n�ԫ��6�1<�D)�$>6��Ds�7P��g�y�R,\n��WA���U��n"0��&���9�_�¸�GSd��U��t���0�0:"�it�Ɇ��;½���[$��k	�&�{�F�����m��iR9U2).����j���T:Ye�X��i̱���k���]�;3�J�Y�z$��%C����4=J�^��Wa���x`5���AVt�U�h�����=����I�o���Gx�6,��o��f��̪�v�W:m�k�>��������Z��]�,b�0��25 �rh�"�/�t���>����%�ѭ�0�.EN� �{[j:�_��b]�����ez&�#]�M����K�f/� 8���"*��1,�g��T��G��u���˙�ބ�_�<�%[|w�&b:F�U����� nȄH���L�ݍ{4J��ڃ�ĺ�;#�o�� e���{��pu@.6��}7݃0_�K6��*<N�����Q��fζҟ|%V��~7V�=|������$���(�o�J����F�d�z�\���rM�x�G�XHb��.��)쌘'׀�0���uN��y�$���+�@�?��#�{�+��ܒ� �t��~��N����@7�1�������S`�?v<��X�o/�ˍ�?Ǯ=��YzPJ��A8�@�����@��,�V��/�;&wP���%�m56W�#����~΄InO�IFW��i!?*�P��&eD݃/�n�D\��&œd�T,�xi��h@��`��9WP���|F�3^�O+O�&��f��
�~	�/���G�9���9+n��L 1��-�}��i?��IҭOQ�2��bpjľ�FM�N.�rr�#��&j#92��$���c���T���������l�S%3�-�#(��У^c6��رܷ��wbP�G�V����~r��$���
b&J���0i:�I�.���a͘=�2��6x����d{�3kҼ��ȼ5����uD��?|&F�%c�O�J�>�˅� �;qW�v��^�!]��e�Ic��J����`-�_uu
��?�gJJ�?�9a!�K�a����F]��G�фb��]rN�wJ�RQ��Ǆt�C��UJ����uI-�A5���|����D��\�H��.�t�7y��$�C�&W�,�x�	Y��B�A�w)�W�R����*I�����c��<G��u�f|m�2-~���73���?��{����N9]�����D�\��:xÎJ&���j�H�%��0NaQ�%�>�^��Z 4�RT����Xj:�ƮB�8+��J�@����,�R$����'bD����4�,'��dDҚy��QX�OcUa�";X��&���Fc˓��� �}|C�> %)�Y2�W��e�h,���ϡ���1m��^�pNu���N(���(�.ŵ�#4��pC��WO�*O�����>&���H��+�/i��Cz�eO�hm���d���>��w2��;��s����[��lE��c�4�Z��Y+��.���!���_�m�g���
d7��V�~�E�0���߂A���L��&�O@m
��9�����{sz�FQ��kKL&˸z��M̦�PM|��c��%~_�
>�oY6�!�,c�Sr���I��2?�Bxl{(Yƀ?�5��򥐿}Z���Pf���Ŕ��Vf�g<�!P؛� ꂙX����/��h��l��_�s>�H.`U6�{��`?��!HT ��^_a��8�G������,�x|=Lq�'cA������z8����4�/�،�e�d��2�=���Ѽ�]h�UvN���iބo�o/��?��Fhe8Tcy���lp=���a����Ɉ\R�Q�p^PveT�9^ٯ�=�3�q?ݢ
���T�4�iT;Cy��6�b�F���F�!���m�K�ۑ2�I���㙤�|S��[��r���a(��1��J*�ȧׯ8�g�;͏pJ��n���'�Du[�
l&�@f�(�"8�ј��5�?_q�ر��n�G��?Ci ���E/�����̬�9��d�+k��w��zs��П�Р��:	Q��W�|���o�!@)�'�, +�vk.�9�j�S� ���}��M�3i�qLA�Y�7��P27X���J0>��s4.�>���"��i�/�`Z��-[��+X�+�w�h�+Ĩ��)A���eqֽ|�6�ܰ�/K��Ro��q*׮�n���cq>T�m&Hu`����?�/%��|�ǜ#��n6�J{�٭��T�D��m���j'���D�r,�1+7�&��'�@iO �yJ���p!{!���{����,0A�C�M���B��81���#��檊� �EH�}G)�� ap�z��l��}�1ρ������ |B|�	��kej+cc�;/� ��*�3㖻 ������%{�H���2	~`�2��a�o�y{�h>W�d�Ls�G�5�����j�Va���{.	�d1	�lT��n�HZ�?��Ӛ�j����w�3��g"Is�U�4�O@s(�Q����zP)fæ
Z� >]%��˼����x�h@<fdp��0�����K � ���/�8~�<Ga��p����a9=�Av�ӚI!�.y\�M\�LZZ���n����	�Jj��r<�E���_�Mp�A�Q�Ck���4t�u�!9>t��:*C2�f��_��ժNOV����WA�.'t�O��N��H{��6+r�ib*b�Gʮ̀�d���誸�(/ǭ��vS�qL�4��9A4��H���<H%,�E]��Z���%�|�K��|�<�Si�U'���4��D+,�G{D�!ke(����gV#]���i���)BjK3RRz�a��hM%j0��e�c{�1�C�<��!���K��������_:��i郤D�*9d��״��G��@�K%�	���ۭ��4�n���*/a��N���/|k�������"��qv:k������޵�#�}{_{�Q�����k���8Y\:\f��Uo���M��,Q77ѐ{��>\\[?�����Q*�3>aO������U:�Ʊ����>Qb�������]U�p����?5������xw�o�7G�'&�r�J�!���)�j�p��:	(�������z,����-�ynm���3H*�o4[�ՙ��&���������eV�	��d����%0=���n,q��j�(�-��� �K|( =f������ {� zR���6L] ��7|>b�N�OB����R�wB����#�Z%�m�2�ɾ1NA�}���t�O�[���T�%Ja{���}dı:�%���8���IO�����Kiw[:��9�`�U����k%�(EJj�^dp�;Y؆�sN�ǶD� ��i�����1g�VG#�-7)�޽9w҂�������h��56˓��BWV�y,M	p�5����9��X��$5��倕D�[�ܚȽ~���TyGx8�q;��}�t��N�� '&=�� ��)QgIwU��	�����Q/m�ҨV#c.����_�����˴~�n䌯Q@�G%��X��`�L�%����O� ��2��k\+vo�����˞�A ��i�Q^�:��r��6���3m�*Ɲ��T�7C:@��I45:�w�X\Q2���t�r
�>����z�-��)tF���W����Bb��$�Yf<]��y���k��\��
�4�`~�}�T��[���"
(�|I�2E���W+�Vtr!c`�9